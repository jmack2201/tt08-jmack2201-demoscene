module sprite_rom1 (
	input clk,
	input [11:0] addr,
	output reg [5:0] color_out
);
	reg [5:0] color_arr [SPRITE_SIZE*SPRITE_SIZE-1:0];

	initial begin
		color_arr[0] = 6'b000000;
		color_arr[1] = 6'b000000;
		color_arr[2] = 6'b000000;
		color_arr[3] = 6'b000000;
		color_arr[4] = 6'b000000;
		color_arr[5] = 6'b000000;
		color_arr[6] = 6'b000000;
		color_arr[7] = 6'b000000;
		color_arr[8] = 6'b000000;
		color_arr[9] = 6'b000000;
		color_arr[10] = 6'b000000;
		color_arr[11] = 6'b000000;
		color_arr[12] = 6'b000000;
		color_arr[13] = 6'b000000;
		color_arr[14] = 6'b000000;
		color_arr[15] = 6'b000000;
		color_arr[16] = 6'b000000;
		color_arr[17] = 6'b000000;
		color_arr[18] = 6'b000000;
		color_arr[19] = 6'b000000;
		color_arr[20] = 6'b000000;
		color_arr[21] = 6'b000000;
		color_arr[22] = 6'b000000;
		color_arr[23] = 6'b000000;
		color_arr[24] = 6'b000000;
		color_arr[25] = 6'b000000;
		color_arr[26] = 6'b000000;
		color_arr[27] = 6'b000000;
		color_arr[28] = 6'b000000;
		color_arr[29] = 6'b000000;
		color_arr[30] = 6'b000000;
		color_arr[31] = 6'b000000;
		color_arr[32] = 6'b000000;
		color_arr[33] = 6'b000000;
		color_arr[34] = 6'b000000;
		color_arr[35] = 6'b000000;
		color_arr[36] = 6'b000000;
		color_arr[37] = 6'b000000;
		color_arr[38] = 6'b000000;
		color_arr[39] = 6'b000000;
		color_arr[40] = 6'b000000;
		color_arr[41] = 6'b000000;
		color_arr[42] = 6'b000000;
		color_arr[43] = 6'b000000;
		color_arr[44] = 6'b000000;
		color_arr[45] = 6'b000000;
		color_arr[46] = 6'b000000;
		color_arr[47] = 6'b000000;
		color_arr[48] = 6'b000000;
		color_arr[49] = 6'b000000;
		color_arr[50] = 6'b000000;
		color_arr[51] = 6'b000000;
		color_arr[52] = 6'b000000;
		color_arr[53] = 6'b000000;
		color_arr[54] = 6'b000000;
		color_arr[55] = 6'b000000;
		color_arr[56] = 6'b000000;
		color_arr[57] = 6'b000000;
		color_arr[58] = 6'b000000;
		color_arr[59] = 6'b000000;
		color_arr[60] = 6'b000000;
		color_arr[61] = 6'b000000;
		color_arr[62] = 6'b000000;
		color_arr[63] = 6'b000000;
		color_arr[64] = 6'b000000;
		color_arr[65] = 6'b000000;
		color_arr[66] = 6'b000000;
		color_arr[67] = 6'b000000;
		color_arr[68] = 6'b000000;
		color_arr[69] = 6'b000000;
		color_arr[70] = 6'b000000;
		color_arr[71] = 6'b000000;
		color_arr[72] = 6'b000000;
		color_arr[73] = 6'b000000;
		color_arr[74] = 6'b000000;
		color_arr[75] = 6'b000000;
		color_arr[76] = 6'b000000;
		color_arr[77] = 6'b000000;
		color_arr[78] = 6'b000000;
		color_arr[79] = 6'b000000;
		color_arr[80] = 6'b000000;
		color_arr[81] = 6'b000000;
		color_arr[82] = 6'b000000;
		color_arr[83] = 6'b000000;
		color_arr[84] = 6'b000000;
		color_arr[85] = 6'b000000;
		color_arr[86] = 6'b000000;
		color_arr[87] = 6'b000000;
		color_arr[88] = 6'b000000;
		color_arr[89] = 6'b000000;
		color_arr[90] = 6'b000000;
		color_arr[91] = 6'b000000;
		color_arr[92] = 6'b000000;
		color_arr[93] = 6'b000000;
		color_arr[94] = 6'b000000;
		color_arr[95] = 6'b000000;
		color_arr[96] = 6'b000000;
		color_arr[97] = 6'b000000;
		color_arr[98] = 6'b000000;
		color_arr[99] = 6'b000000;
		color_arr[100] = 6'b000000;
		color_arr[101] = 6'b000000;
		color_arr[102] = 6'b000000;
		color_arr[103] = 6'b000000;
		color_arr[104] = 6'b000000;
		color_arr[105] = 6'b000000;
		color_arr[106] = 6'b000000;
		color_arr[107] = 6'b000000;
		color_arr[108] = 6'b000000;
		color_arr[109] = 6'b000000;
		color_arr[110] = 6'b000000;
		color_arr[111] = 6'b000000;
		color_arr[112] = 6'b000000;
		color_arr[113] = 6'b000000;
		color_arr[114] = 6'b000000;
		color_arr[115] = 6'b000000;
		color_arr[116] = 6'b000000;
		color_arr[117] = 6'b000000;
		color_arr[118] = 6'b000000;
		color_arr[119] = 6'b000000;
		color_arr[120] = 6'b000000;
		color_arr[121] = 6'b000000;
		color_arr[122] = 6'b000000;
		color_arr[123] = 6'b000000;
		color_arr[124] = 6'b000000;
		color_arr[125] = 6'b000000;
		color_arr[126] = 6'b000000;
		color_arr[127] = 6'b000000;
		color_arr[128] = 6'b000000;
		color_arr[129] = 6'b000000;
		color_arr[130] = 6'b000000;
		color_arr[131] = 6'b000000;
		color_arr[132] = 6'b000000;
		color_arr[133] = 6'b000000;
		color_arr[134] = 6'b000000;
		color_arr[135] = 6'b000000;
		color_arr[136] = 6'b000000;
		color_arr[137] = 6'b000000;
		color_arr[138] = 6'b000000;
		color_arr[139] = 6'b000000;
		color_arr[140] = 6'b000000;
		color_arr[141] = 6'b000000;
		color_arr[142] = 6'b000000;
		color_arr[143] = 6'b000000;
		color_arr[144] = 6'b000000;
		color_arr[145] = 6'b000000;
		color_arr[146] = 6'b000000;
		color_arr[147] = 6'b000000;
		color_arr[148] = 6'b000000;
		color_arr[149] = 6'b000000;
		color_arr[150] = 6'b000000;
		color_arr[151] = 6'b000000;
		color_arr[152] = 6'b000000;
		color_arr[153] = 6'b000000;
		color_arr[154] = 6'b000000;
		color_arr[155] = 6'b000000;
		color_arr[156] = 6'b000000;
		color_arr[157] = 6'b000000;
		color_arr[158] = 6'b000000;
		color_arr[159] = 6'b000000;
		color_arr[160] = 6'b000000;
		color_arr[161] = 6'b000000;
		color_arr[162] = 6'b000000;
		color_arr[163] = 6'b000000;
		color_arr[164] = 6'b000000;
		color_arr[165] = 6'b000000;
		color_arr[166] = 6'b000000;
		color_arr[167] = 6'b000000;
		color_arr[168] = 6'b000000;
		color_arr[169] = 6'b000000;
		color_arr[170] = 6'b000000;
		color_arr[171] = 6'b000000;
		color_arr[172] = 6'b000000;
		color_arr[173] = 6'b000000;
		color_arr[174] = 6'b000000;
		color_arr[175] = 6'b000000;
		color_arr[176] = 6'b000000;
		color_arr[177] = 6'b000000;
		color_arr[178] = 6'b000000;
		color_arr[179] = 6'b000000;
		color_arr[180] = 6'b000000;
		color_arr[181] = 6'b000000;
		color_arr[182] = 6'b000000;
		color_arr[183] = 6'b000000;
		color_arr[184] = 6'b000000;
		color_arr[185] = 6'b000000;
		color_arr[186] = 6'b000000;
		color_arr[187] = 6'b000000;
		color_arr[188] = 6'b000000;
		color_arr[189] = 6'b000000;
		color_arr[190] = 6'b000000;
		color_arr[191] = 6'b000000;
		color_arr[192] = 6'b000000;
		color_arr[193] = 6'b000000;
		color_arr[194] = 6'b000000;
		color_arr[195] = 6'b000000;
		color_arr[196] = 6'b000000;
		color_arr[197] = 6'b000000;
		color_arr[198] = 6'b000000;
		color_arr[199] = 6'b000000;
		color_arr[200] = 6'b000000;
		color_arr[201] = 6'b000000;
		color_arr[202] = 6'b000000;
		color_arr[203] = 6'b000000;
		color_arr[204] = 6'b000000;
		color_arr[205] = 6'b000000;
		color_arr[206] = 6'b000000;
		color_arr[207] = 6'b000000;
		color_arr[208] = 6'b000000;
		color_arr[209] = 6'b000000;
		color_arr[210] = 6'b000000;
		color_arr[211] = 6'b000000;
		color_arr[212] = 6'b000000;
		color_arr[213] = 6'b000000;
		color_arr[214] = 6'b000000;
		color_arr[215] = 6'b000000;
		color_arr[216] = 6'b000000;
		color_arr[217] = 6'b000000;
		color_arr[218] = 6'b000000;
		color_arr[219] = 6'b000000;
		color_arr[220] = 6'b000000;
		color_arr[221] = 6'b000000;
		color_arr[222] = 6'b000000;
		color_arr[223] = 6'b000000;
		color_arr[224] = 6'b000000;
		color_arr[225] = 6'b000000;
		color_arr[226] = 6'b000000;
		color_arr[227] = 6'b000000;
		color_arr[228] = 6'b000000;
		color_arr[229] = 6'b000000;
		color_arr[230] = 6'b000000;
		color_arr[231] = 6'b000000;
		color_arr[232] = 6'b000000;
		color_arr[233] = 6'b000000;
		color_arr[234] = 6'b000000;
		color_arr[235] = 6'b000000;
		color_arr[236] = 6'b000000;
		color_arr[237] = 6'b000000;
		color_arr[238] = 6'b000000;
		color_arr[239] = 6'b000000;
		color_arr[240] = 6'b000000;
		color_arr[241] = 6'b000000;
		color_arr[242] = 6'b000000;
		color_arr[243] = 6'b000000;
		color_arr[244] = 6'b000000;
		color_arr[245] = 6'b000000;
		color_arr[246] = 6'b000000;
		color_arr[247] = 6'b000000;
		color_arr[248] = 6'b000000;
		color_arr[249] = 6'b000000;
		color_arr[250] = 6'b000000;
		color_arr[251] = 6'b000000;
		color_arr[252] = 6'b000000;
		color_arr[253] = 6'b000000;
		color_arr[254] = 6'b000000;
		color_arr[255] = 6'b000000;
		color_arr[256] = 6'b000000;
		color_arr[257] = 6'b000000;
		color_arr[258] = 6'b000000;
		color_arr[259] = 6'b000000;
		color_arr[260] = 6'b000000;
		color_arr[261] = 6'b000000;
		color_arr[262] = 6'b000000;
		color_arr[263] = 6'b000000;
		color_arr[264] = 6'b000000;
		color_arr[265] = 6'b000000;
		color_arr[266] = 6'b000000;
		color_arr[267] = 6'b000000;
		color_arr[268] = 6'b000000;
		color_arr[269] = 6'b000000;
		color_arr[270] = 6'b000000;
		color_arr[271] = 6'b000000;
		color_arr[272] = 6'b000000;
		color_arr[273] = 6'b000000;
		color_arr[274] = 6'b000000;
		color_arr[275] = 6'b000000;
		color_arr[276] = 6'b000000;
		color_arr[277] = 6'b000000;
		color_arr[278] = 6'b000000;
		color_arr[279] = 6'b000000;
		color_arr[280] = 6'b000000;
		color_arr[281] = 6'b000000;
		color_arr[282] = 6'b000000;
		color_arr[283] = 6'b000000;
		color_arr[284] = 6'b000000;
		color_arr[285] = 6'b000000;
		color_arr[286] = 6'b000000;
		color_arr[287] = 6'b000000;
		color_arr[288] = 6'b000000;
		color_arr[289] = 6'b000000;
		color_arr[290] = 6'b000000;
		color_arr[291] = 6'b000000;
		color_arr[292] = 6'b000000;
		color_arr[293] = 6'b000000;
		color_arr[294] = 6'b000000;
		color_arr[295] = 6'b000000;
		color_arr[296] = 6'b000000;
		color_arr[297] = 6'b000000;
		color_arr[298] = 6'b000000;
		color_arr[299] = 6'b000000;
		color_arr[300] = 6'b000000;
		color_arr[301] = 6'b000000;
		color_arr[302] = 6'b000000;
		color_arr[303] = 6'b000000;
		color_arr[304] = 6'b000000;
		color_arr[305] = 6'b000000;
		color_arr[306] = 6'b000000;
		color_arr[307] = 6'b000000;
		color_arr[308] = 6'b000000;
		color_arr[309] = 6'b000000;
		color_arr[310] = 6'b000000;
		color_arr[311] = 6'b000000;
		color_arr[312] = 6'b000000;
		color_arr[313] = 6'b000000;
		color_arr[314] = 6'b000000;
		color_arr[315] = 6'b000000;
		color_arr[316] = 6'b000000;
		color_arr[317] = 6'b000000;
		color_arr[318] = 6'b000000;
		color_arr[319] = 6'b000000;
		color_arr[320] = 6'b000000;
		color_arr[321] = 6'b000000;
		color_arr[322] = 6'b000000;
		color_arr[323] = 6'b000000;
		color_arr[324] = 6'b000000;
		color_arr[325] = 6'b000000;
		color_arr[326] = 6'b000000;
		color_arr[327] = 6'b000000;
		color_arr[328] = 6'b000000;
		color_arr[329] = 6'b000000;
		color_arr[330] = 6'b000000;
		color_arr[331] = 6'b000000;
		color_arr[332] = 6'b000000;
		color_arr[333] = 6'b000000;
		color_arr[334] = 6'b000000;
		color_arr[335] = 6'b000000;
		color_arr[336] = 6'b000000;
		color_arr[337] = 6'b000000;
		color_arr[338] = 6'b000000;
		color_arr[339] = 6'b000000;
		color_arr[340] = 6'b000000;
		color_arr[341] = 6'b000000;
		color_arr[342] = 6'b111001;
		color_arr[343] = 6'b000000;
		color_arr[344] = 6'b000000;
		color_arr[345] = 6'b000000;
		color_arr[346] = 6'b000000;
		color_arr[347] = 6'b000000;
		color_arr[348] = 6'b000000;
		color_arr[349] = 6'b000000;
		color_arr[350] = 6'b000000;
		color_arr[351] = 6'b000000;
		color_arr[352] = 6'b000000;
		color_arr[353] = 6'b000000;
		color_arr[354] = 6'b000000;
		color_arr[355] = 6'b000000;
		color_arr[356] = 6'b000000;
		color_arr[357] = 6'b000000;
		color_arr[358] = 6'b000000;
		color_arr[359] = 6'b000000;
		color_arr[360] = 6'b000000;
		color_arr[361] = 6'b000000;
		color_arr[362] = 6'b000000;
		color_arr[363] = 6'b000000;
		color_arr[364] = 6'b000000;
		color_arr[365] = 6'b000000;
		color_arr[366] = 6'b000000;
		color_arr[367] = 6'b000000;
		color_arr[368] = 6'b000000;
		color_arr[369] = 6'b000000;
		color_arr[370] = 6'b000000;
		color_arr[371] = 6'b000000;
		color_arr[372] = 6'b000000;
		color_arr[373] = 6'b000000;
		color_arr[374] = 6'b000000;
		color_arr[375] = 6'b000000;
		color_arr[376] = 6'b000000;
		color_arr[377] = 6'b000000;
		color_arr[378] = 6'b000000;
		color_arr[379] = 6'b000000;
		color_arr[380] = 6'b000000;
		color_arr[381] = 6'b000000;
		color_arr[382] = 6'b000000;
		color_arr[383] = 6'b000000;
		color_arr[384] = 6'b000000;
		color_arr[385] = 6'b000000;
		color_arr[386] = 6'b000000;
		color_arr[387] = 6'b000000;
		color_arr[388] = 6'b000000;
		color_arr[389] = 6'b000000;
		color_arr[390] = 6'b000000;
		color_arr[391] = 6'b000000;
		color_arr[392] = 6'b000000;
		color_arr[393] = 6'b000000;
		color_arr[394] = 6'b000000;
		color_arr[395] = 6'b000000;
		color_arr[396] = 6'b000000;
		color_arr[397] = 6'b000000;
		color_arr[398] = 6'b000000;
		color_arr[399] = 6'b000000;
		color_arr[400] = 6'b000000;
		color_arr[401] = 6'b000000;
		color_arr[402] = 6'b000000;
		color_arr[403] = 6'b000000;
		color_arr[404] = 6'b000000;
		color_arr[405] = 6'b101000;
		color_arr[406] = 6'b111001;
		color_arr[407] = 6'b111001;
		color_arr[408] = 6'b000000;
		color_arr[409] = 6'b000000;
		color_arr[410] = 6'b000000;
		color_arr[411] = 6'b000000;
		color_arr[412] = 6'b000000;
		color_arr[413] = 6'b000000;
		color_arr[414] = 6'b000000;
		color_arr[415] = 6'b000000;
		color_arr[416] = 6'b000000;
		color_arr[417] = 6'b000000;
		color_arr[418] = 6'b000000;
		color_arr[419] = 6'b000000;
		color_arr[420] = 6'b111001;
		color_arr[421] = 6'b000000;
		color_arr[422] = 6'b000000;
		color_arr[423] = 6'b000000;
		color_arr[424] = 6'b000000;
		color_arr[425] = 6'b000000;
		color_arr[426] = 6'b000000;
		color_arr[427] = 6'b000000;
		color_arr[428] = 6'b000000;
		color_arr[429] = 6'b000000;
		color_arr[430] = 6'b000000;
		color_arr[431] = 6'b000000;
		color_arr[432] = 6'b000000;
		color_arr[433] = 6'b000000;
		color_arr[434] = 6'b000000;
		color_arr[435] = 6'b000000;
		color_arr[436] = 6'b000000;
		color_arr[437] = 6'b000000;
		color_arr[438] = 6'b000000;
		color_arr[439] = 6'b000000;
		color_arr[440] = 6'b000000;
		color_arr[441] = 6'b000000;
		color_arr[442] = 6'b000000;
		color_arr[443] = 6'b000000;
		color_arr[444] = 6'b000000;
		color_arr[445] = 6'b000000;
		color_arr[446] = 6'b000000;
		color_arr[447] = 6'b000000;
		color_arr[448] = 6'b000000;
		color_arr[449] = 6'b000000;
		color_arr[450] = 6'b000000;
		color_arr[451] = 6'b000000;
		color_arr[452] = 6'b000000;
		color_arr[453] = 6'b000000;
		color_arr[454] = 6'b000000;
		color_arr[455] = 6'b000000;
		color_arr[456] = 6'b000000;
		color_arr[457] = 6'b000000;
		color_arr[458] = 6'b000000;
		color_arr[459] = 6'b000000;
		color_arr[460] = 6'b000000;
		color_arr[461] = 6'b000000;
		color_arr[462] = 6'b000000;
		color_arr[463] = 6'b000000;
		color_arr[464] = 6'b000000;
		color_arr[465] = 6'b000000;
		color_arr[466] = 6'b000000;
		color_arr[467] = 6'b000000;
		color_arr[468] = 6'b000000;
		color_arr[469] = 6'b101000;
		color_arr[470] = 6'b111001;
		color_arr[471] = 6'b111001;
		color_arr[472] = 6'b000000;
		color_arr[473] = 6'b000000;
		color_arr[474] = 6'b000000;
		color_arr[475] = 6'b000000;
		color_arr[476] = 6'b000000;
		color_arr[477] = 6'b000000;
		color_arr[478] = 6'b000000;
		color_arr[479] = 6'b000000;
		color_arr[480] = 6'b000000;
		color_arr[481] = 6'b000000;
		color_arr[482] = 6'b000000;
		color_arr[483] = 6'b111001;
		color_arr[484] = 6'b111001;
		color_arr[485] = 6'b111001;
		color_arr[486] = 6'b000000;
		color_arr[487] = 6'b000000;
		color_arr[488] = 6'b000000;
		color_arr[489] = 6'b000000;
		color_arr[490] = 6'b000000;
		color_arr[491] = 6'b000000;
		color_arr[492] = 6'b000000;
		color_arr[493] = 6'b000000;
		color_arr[494] = 6'b000000;
		color_arr[495] = 6'b000000;
		color_arr[496] = 6'b000000;
		color_arr[497] = 6'b000000;
		color_arr[498] = 6'b000000;
		color_arr[499] = 6'b000000;
		color_arr[500] = 6'b000000;
		color_arr[501] = 6'b000000;
		color_arr[502] = 6'b000000;
		color_arr[503] = 6'b000000;
		color_arr[504] = 6'b000000;
		color_arr[505] = 6'b000000;
		color_arr[506] = 6'b000000;
		color_arr[507] = 6'b000000;
		color_arr[508] = 6'b000000;
		color_arr[509] = 6'b000000;
		color_arr[510] = 6'b000000;
		color_arr[511] = 6'b000000;
		color_arr[512] = 6'b000000;
		color_arr[513] = 6'b000000;
		color_arr[514] = 6'b000000;
		color_arr[515] = 6'b000000;
		color_arr[516] = 6'b000000;
		color_arr[517] = 6'b000000;
		color_arr[518] = 6'b000000;
		color_arr[519] = 6'b000000;
		color_arr[520] = 6'b000000;
		color_arr[521] = 6'b000000;
		color_arr[522] = 6'b000000;
		color_arr[523] = 6'b000000;
		color_arr[524] = 6'b000000;
		color_arr[525] = 6'b000000;
		color_arr[526] = 6'b000000;
		color_arr[527] = 6'b000000;
		color_arr[528] = 6'b000000;
		color_arr[529] = 6'b000000;
		color_arr[530] = 6'b000000;
		color_arr[531] = 6'b000000;
		color_arr[532] = 6'b000000;
		color_arr[533] = 6'b101000;
		color_arr[534] = 6'b111001;
		color_arr[535] = 6'b111001;
		color_arr[536] = 6'b111001;
		color_arr[537] = 6'b000000;
		color_arr[538] = 6'b000000;
		color_arr[539] = 6'b000000;
		color_arr[540] = 6'b000000;
		color_arr[541] = 6'b000000;
		color_arr[542] = 6'b000000;
		color_arr[543] = 6'b000000;
		color_arr[544] = 6'b000000;
		color_arr[545] = 6'b000000;
		color_arr[546] = 6'b111001;
		color_arr[547] = 6'b111001;
		color_arr[548] = 6'b111001;
		color_arr[549] = 6'b111001;
		color_arr[550] = 6'b000000;
		color_arr[551] = 6'b000000;
		color_arr[552] = 6'b000000;
		color_arr[553] = 6'b000000;
		color_arr[554] = 6'b000000;
		color_arr[555] = 6'b000000;
		color_arr[556] = 6'b000000;
		color_arr[557] = 6'b000000;
		color_arr[558] = 6'b000000;
		color_arr[559] = 6'b000000;
		color_arr[560] = 6'b000000;
		color_arr[561] = 6'b000000;
		color_arr[562] = 6'b000000;
		color_arr[563] = 6'b000000;
		color_arr[564] = 6'b000000;
		color_arr[565] = 6'b000000;
		color_arr[566] = 6'b000000;
		color_arr[567] = 6'b000000;
		color_arr[568] = 6'b000000;
		color_arr[569] = 6'b000000;
		color_arr[570] = 6'b000000;
		color_arr[571] = 6'b000000;
		color_arr[572] = 6'b000000;
		color_arr[573] = 6'b000000;
		color_arr[574] = 6'b000000;
		color_arr[575] = 6'b000000;
		color_arr[576] = 6'b000000;
		color_arr[577] = 6'b000000;
		color_arr[578] = 6'b000000;
		color_arr[579] = 6'b000000;
		color_arr[580] = 6'b000000;
		color_arr[581] = 6'b000000;
		color_arr[582] = 6'b000000;
		color_arr[583] = 6'b000000;
		color_arr[584] = 6'b000000;
		color_arr[585] = 6'b000000;
		color_arr[586] = 6'b000000;
		color_arr[587] = 6'b000000;
		color_arr[588] = 6'b000000;
		color_arr[589] = 6'b000000;
		color_arr[590] = 6'b000000;
		color_arr[591] = 6'b000000;
		color_arr[592] = 6'b000000;
		color_arr[593] = 6'b000000;
		color_arr[594] = 6'b000000;
		color_arr[595] = 6'b000000;
		color_arr[596] = 6'b000000;
		color_arr[597] = 6'b111001;
		color_arr[598] = 6'b111001;
		color_arr[599] = 6'b111001;
		color_arr[600] = 6'b111001;
		color_arr[601] = 6'b111001;
		color_arr[602] = 6'b111001;
		color_arr[603] = 6'b000000;
		color_arr[604] = 6'b000000;
		color_arr[605] = 6'b000000;
		color_arr[606] = 6'b000000;
		color_arr[607] = 6'b000000;
		color_arr[608] = 6'b111001;
		color_arr[609] = 6'b111001;
		color_arr[610] = 6'b111001;
		color_arr[611] = 6'b111001;
		color_arr[612] = 6'b101000;
		color_arr[613] = 6'b111001;
		color_arr[614] = 6'b111001;
		color_arr[615] = 6'b000000;
		color_arr[616] = 6'b000000;
		color_arr[617] = 6'b000000;
		color_arr[618] = 6'b000000;
		color_arr[619] = 6'b000000;
		color_arr[620] = 6'b000000;
		color_arr[621] = 6'b000000;
		color_arr[622] = 6'b000000;
		color_arr[623] = 6'b000000;
		color_arr[624] = 6'b000000;
		color_arr[625] = 6'b000000;
		color_arr[626] = 6'b000000;
		color_arr[627] = 6'b000000;
		color_arr[628] = 6'b000000;
		color_arr[629] = 6'b000000;
		color_arr[630] = 6'b000000;
		color_arr[631] = 6'b000000;
		color_arr[632] = 6'b000000;
		color_arr[633] = 6'b000000;
		color_arr[634] = 6'b000000;
		color_arr[635] = 6'b000000;
		color_arr[636] = 6'b000000;
		color_arr[637] = 6'b000000;
		color_arr[638] = 6'b000000;
		color_arr[639] = 6'b000000;
		color_arr[640] = 6'b000000;
		color_arr[641] = 6'b000000;
		color_arr[642] = 6'b000000;
		color_arr[643] = 6'b000000;
		color_arr[644] = 6'b000000;
		color_arr[645] = 6'b000000;
		color_arr[646] = 6'b000000;
		color_arr[647] = 6'b000000;
		color_arr[648] = 6'b000000;
		color_arr[649] = 6'b000000;
		color_arr[650] = 6'b000000;
		color_arr[651] = 6'b000000;
		color_arr[652] = 6'b000000;
		color_arr[653] = 6'b000000;
		color_arr[654] = 6'b000000;
		color_arr[655] = 6'b000000;
		color_arr[656] = 6'b000000;
		color_arr[657] = 6'b000000;
		color_arr[658] = 6'b000000;
		color_arr[659] = 6'b000000;
		color_arr[660] = 6'b111001;
		color_arr[661] = 6'b111001;
		color_arr[662] = 6'b111001;
		color_arr[663] = 6'b111001;
		color_arr[664] = 6'b111001;
		color_arr[665] = 6'b111001;
		color_arr[666] = 6'b111001;
		color_arr[667] = 6'b111001;
		color_arr[668] = 6'b111001;
		color_arr[669] = 6'b111001;
		color_arr[670] = 6'b111001;
		color_arr[671] = 6'b111001;
		color_arr[672] = 6'b111001;
		color_arr[673] = 6'b111001;
		color_arr[674] = 6'b111001;
		color_arr[675] = 6'b111001;
		color_arr[676] = 6'b101000;
		color_arr[677] = 6'b111001;
		color_arr[678] = 6'b111001;
		color_arr[679] = 6'b111001;
		color_arr[680] = 6'b000000;
		color_arr[681] = 6'b000000;
		color_arr[682] = 6'b000000;
		color_arr[683] = 6'b000000;
		color_arr[684] = 6'b000000;
		color_arr[685] = 6'b000000;
		color_arr[686] = 6'b000000;
		color_arr[687] = 6'b000000;
		color_arr[688] = 6'b000000;
		color_arr[689] = 6'b000000;
		color_arr[690] = 6'b000000;
		color_arr[691] = 6'b000000;
		color_arr[692] = 6'b000000;
		color_arr[693] = 6'b000000;
		color_arr[694] = 6'b000000;
		color_arr[695] = 6'b000000;
		color_arr[696] = 6'b000000;
		color_arr[697] = 6'b000000;
		color_arr[698] = 6'b000000;
		color_arr[699] = 6'b000000;
		color_arr[700] = 6'b000000;
		color_arr[701] = 6'b000000;
		color_arr[702] = 6'b000000;
		color_arr[703] = 6'b000000;
		color_arr[704] = 6'b000000;
		color_arr[705] = 6'b000000;
		color_arr[706] = 6'b000000;
		color_arr[707] = 6'b000000;
		color_arr[708] = 6'b000000;
		color_arr[709] = 6'b000000;
		color_arr[710] = 6'b000000;
		color_arr[711] = 6'b000000;
		color_arr[712] = 6'b000000;
		color_arr[713] = 6'b000000;
		color_arr[714] = 6'b000000;
		color_arr[715] = 6'b000000;
		color_arr[716] = 6'b000000;
		color_arr[717] = 6'b000000;
		color_arr[718] = 6'b000000;
		color_arr[719] = 6'b000000;
		color_arr[720] = 6'b000000;
		color_arr[721] = 6'b000000;
		color_arr[722] = 6'b000000;
		color_arr[723] = 6'b111001;
		color_arr[724] = 6'b111001;
		color_arr[725] = 6'b111001;
		color_arr[726] = 6'b111001;
		color_arr[727] = 6'b111001;
		color_arr[728] = 6'b111001;
		color_arr[729] = 6'b111001;
		color_arr[730] = 6'b111001;
		color_arr[731] = 6'b111001;
		color_arr[732] = 6'b111001;
		color_arr[733] = 6'b111001;
		color_arr[734] = 6'b111001;
		color_arr[735] = 6'b111001;
		color_arr[736] = 6'b111001;
		color_arr[737] = 6'b111001;
		color_arr[738] = 6'b111001;
		color_arr[739] = 6'b101000;
		color_arr[740] = 6'b101000;
		color_arr[741] = 6'b111001;
		color_arr[742] = 6'b111001;
		color_arr[743] = 6'b111001;
		color_arr[744] = 6'b000000;
		color_arr[745] = 6'b000000;
		color_arr[746] = 6'b000000;
		color_arr[747] = 6'b000000;
		color_arr[748] = 6'b000000;
		color_arr[749] = 6'b000000;
		color_arr[750] = 6'b000000;
		color_arr[751] = 6'b000000;
		color_arr[752] = 6'b000000;
		color_arr[753] = 6'b000000;
		color_arr[754] = 6'b000000;
		color_arr[755] = 6'b000000;
		color_arr[756] = 6'b000000;
		color_arr[757] = 6'b000000;
		color_arr[758] = 6'b000000;
		color_arr[759] = 6'b000000;
		color_arr[760] = 6'b000000;
		color_arr[761] = 6'b000000;
		color_arr[762] = 6'b000000;
		color_arr[763] = 6'b000000;
		color_arr[764] = 6'b000000;
		color_arr[765] = 6'b000000;
		color_arr[766] = 6'b000000;
		color_arr[767] = 6'b000000;
		color_arr[768] = 6'b000000;
		color_arr[769] = 6'b000000;
		color_arr[770] = 6'b000000;
		color_arr[771] = 6'b000000;
		color_arr[772] = 6'b000000;
		color_arr[773] = 6'b000000;
		color_arr[774] = 6'b000000;
		color_arr[775] = 6'b000000;
		color_arr[776] = 6'b000000;
		color_arr[777] = 6'b000000;
		color_arr[778] = 6'b000000;
		color_arr[779] = 6'b000000;
		color_arr[780] = 6'b000000;
		color_arr[781] = 6'b000000;
		color_arr[782] = 6'b000000;
		color_arr[783] = 6'b000000;
		color_arr[784] = 6'b000000;
		color_arr[785] = 6'b000000;
		color_arr[786] = 6'b111001;
		color_arr[787] = 6'b111001;
		color_arr[788] = 6'b111001;
		color_arr[789] = 6'b111001;
		color_arr[790] = 6'b111001;
		color_arr[791] = 6'b111110;
		color_arr[792] = 6'b111001;
		color_arr[793] = 6'b111001;
		color_arr[794] = 6'b111001;
		color_arr[795] = 6'b111001;
		color_arr[796] = 6'b111001;
		color_arr[797] = 6'b111001;
		color_arr[798] = 6'b111001;
		color_arr[799] = 6'b111001;
		color_arr[800] = 6'b111001;
		color_arr[801] = 6'b111001;
		color_arr[802] = 6'b111001;
		color_arr[803] = 6'b111001;
		color_arr[804] = 6'b111001;
		color_arr[805] = 6'b111001;
		color_arr[806] = 6'b111001;
		color_arr[807] = 6'b111001;
		color_arr[808] = 6'b111001;
		color_arr[809] = 6'b000000;
		color_arr[810] = 6'b000000;
		color_arr[811] = 6'b000000;
		color_arr[812] = 6'b000000;
		color_arr[813] = 6'b000000;
		color_arr[814] = 6'b000000;
		color_arr[815] = 6'b000000;
		color_arr[816] = 6'b000000;
		color_arr[817] = 6'b000000;
		color_arr[818] = 6'b000000;
		color_arr[819] = 6'b000000;
		color_arr[820] = 6'b000000;
		color_arr[821] = 6'b000000;
		color_arr[822] = 6'b000000;
		color_arr[823] = 6'b000000;
		color_arr[824] = 6'b000000;
		color_arr[825] = 6'b000000;
		color_arr[826] = 6'b000000;
		color_arr[827] = 6'b000000;
		color_arr[828] = 6'b000000;
		color_arr[829] = 6'b000000;
		color_arr[830] = 6'b000000;
		color_arr[831] = 6'b000000;
		color_arr[832] = 6'b000000;
		color_arr[833] = 6'b000000;
		color_arr[834] = 6'b000000;
		color_arr[835] = 6'b000000;
		color_arr[836] = 6'b000000;
		color_arr[837] = 6'b000000;
		color_arr[838] = 6'b000000;
		color_arr[839] = 6'b000000;
		color_arr[840] = 6'b000000;
		color_arr[841] = 6'b000000;
		color_arr[842] = 6'b000000;
		color_arr[843] = 6'b000000;
		color_arr[844] = 6'b000000;
		color_arr[845] = 6'b000000;
		color_arr[846] = 6'b000000;
		color_arr[847] = 6'b000000;
		color_arr[848] = 6'b000000;
		color_arr[849] = 6'b111001;
		color_arr[850] = 6'b111001;
		color_arr[851] = 6'b111001;
		color_arr[852] = 6'b111001;
		color_arr[853] = 6'b111001;
		color_arr[854] = 6'b111111;
		color_arr[855] = 6'b111110;
		color_arr[856] = 6'b111001;
		color_arr[857] = 6'b111001;
		color_arr[858] = 6'b111001;
		color_arr[859] = 6'b111001;
		color_arr[860] = 6'b111001;
		color_arr[861] = 6'b111001;
		color_arr[862] = 6'b111110;
		color_arr[863] = 6'b111001;
		color_arr[864] = 6'b111001;
		color_arr[865] = 6'b111001;
		color_arr[866] = 6'b111001;
		color_arr[867] = 6'b111001;
		color_arr[868] = 6'b111001;
		color_arr[869] = 6'b111001;
		color_arr[870] = 6'b111001;
		color_arr[871] = 6'b111001;
		color_arr[872] = 6'b111001;
		color_arr[873] = 6'b000000;
		color_arr[874] = 6'b000000;
		color_arr[875] = 6'b000000;
		color_arr[876] = 6'b000000;
		color_arr[877] = 6'b000000;
		color_arr[878] = 6'b000000;
		color_arr[879] = 6'b000000;
		color_arr[880] = 6'b000000;
		color_arr[881] = 6'b000000;
		color_arr[882] = 6'b000000;
		color_arr[883] = 6'b000000;
		color_arr[884] = 6'b000000;
		color_arr[885] = 6'b000000;
		color_arr[886] = 6'b000000;
		color_arr[887] = 6'b000000;
		color_arr[888] = 6'b000000;
		color_arr[889] = 6'b000000;
		color_arr[890] = 6'b000000;
		color_arr[891] = 6'b000000;
		color_arr[892] = 6'b000000;
		color_arr[893] = 6'b000000;
		color_arr[894] = 6'b000000;
		color_arr[895] = 6'b000000;
		color_arr[896] = 6'b000000;
		color_arr[897] = 6'b000000;
		color_arr[898] = 6'b000000;
		color_arr[899] = 6'b000000;
		color_arr[900] = 6'b000000;
		color_arr[901] = 6'b000000;
		color_arr[902] = 6'b000000;
		color_arr[903] = 6'b000000;
		color_arr[904] = 6'b000000;
		color_arr[905] = 6'b000000;
		color_arr[906] = 6'b000000;
		color_arr[907] = 6'b000000;
		color_arr[908] = 6'b000000;
		color_arr[909] = 6'b000000;
		color_arr[910] = 6'b000000;
		color_arr[911] = 6'b000000;
		color_arr[912] = 6'b000000;
		color_arr[913] = 6'b111001;
		color_arr[914] = 6'b111001;
		color_arr[915] = 6'b111001;
		color_arr[916] = 6'b111001;
		color_arr[917] = 6'b111111;
		color_arr[918] = 6'b111111;
		color_arr[919] = 6'b111110;
		color_arr[920] = 6'b111001;
		color_arr[921] = 6'b111001;
		color_arr[922] = 6'b111001;
		color_arr[923] = 6'b111001;
		color_arr[924] = 6'b111001;
		color_arr[925] = 6'b111110;
		color_arr[926] = 6'b111110;
		color_arr[927] = 6'b111110;
		color_arr[928] = 6'b111110;
		color_arr[929] = 6'b111001;
		color_arr[930] = 6'b111001;
		color_arr[931] = 6'b111001;
		color_arr[932] = 6'b111001;
		color_arr[933] = 6'b111001;
		color_arr[934] = 6'b111001;
		color_arr[935] = 6'b111001;
		color_arr[936] = 6'b111001;
		color_arr[937] = 6'b000000;
		color_arr[938] = 6'b000000;
		color_arr[939] = 6'b000000;
		color_arr[940] = 6'b000000;
		color_arr[941] = 6'b000000;
		color_arr[942] = 6'b000000;
		color_arr[943] = 6'b000000;
		color_arr[944] = 6'b000000;
		color_arr[945] = 6'b000000;
		color_arr[946] = 6'b000000;
		color_arr[947] = 6'b000000;
		color_arr[948] = 6'b000000;
		color_arr[949] = 6'b000000;
		color_arr[950] = 6'b000000;
		color_arr[951] = 6'b000000;
		color_arr[952] = 6'b000000;
		color_arr[953] = 6'b000000;
		color_arr[954] = 6'b000000;
		color_arr[955] = 6'b000000;
		color_arr[956] = 6'b000000;
		color_arr[957] = 6'b000000;
		color_arr[958] = 6'b000000;
		color_arr[959] = 6'b000000;
		color_arr[960] = 6'b000000;
		color_arr[961] = 6'b000000;
		color_arr[962] = 6'b000000;
		color_arr[963] = 6'b000000;
		color_arr[964] = 6'b000000;
		color_arr[965] = 6'b000000;
		color_arr[966] = 6'b000000;
		color_arr[967] = 6'b000000;
		color_arr[968] = 6'b000000;
		color_arr[969] = 6'b000000;
		color_arr[970] = 6'b000000;
		color_arr[971] = 6'b000000;
		color_arr[972] = 6'b000000;
		color_arr[973] = 6'b000000;
		color_arr[974] = 6'b000000;
		color_arr[975] = 6'b000000;
		color_arr[976] = 6'b111001;
		color_arr[977] = 6'b111001;
		color_arr[978] = 6'b111001;
		color_arr[979] = 6'b111001;
		color_arr[980] = 6'b111110;
		color_arr[981] = 6'b111111;
		color_arr[982] = 6'b000000;
		color_arr[983] = 6'b111110;
		color_arr[984] = 6'b111001;
		color_arr[985] = 6'b111001;
		color_arr[986] = 6'b111001;
		color_arr[987] = 6'b111001;
		color_arr[988] = 6'b111001;
		color_arr[989] = 6'b111111;
		color_arr[990] = 6'b111111;
		color_arr[991] = 6'b111111;
		color_arr[992] = 6'b111110;
		color_arr[993] = 6'b111010;
		color_arr[994] = 6'b111010;
		color_arr[995] = 6'b111010;
		color_arr[996] = 6'b111010;
		color_arr[997] = 6'b111001;
		color_arr[998] = 6'b111001;
		color_arr[999] = 6'b111001;
		color_arr[1000] = 6'b111001;
		color_arr[1001] = 6'b000000;
		color_arr[1002] = 6'b000000;
		color_arr[1003] = 6'b000000;
		color_arr[1004] = 6'b000000;
		color_arr[1005] = 6'b000000;
		color_arr[1006] = 6'b000000;
		color_arr[1007] = 6'b000000;
		color_arr[1008] = 6'b000000;
		color_arr[1009] = 6'b000000;
		color_arr[1010] = 6'b000000;
		color_arr[1011] = 6'b000000;
		color_arr[1012] = 6'b000000;
		color_arr[1013] = 6'b000000;
		color_arr[1014] = 6'b000000;
		color_arr[1015] = 6'b000000;
		color_arr[1016] = 6'b000000;
		color_arr[1017] = 6'b000000;
		color_arr[1018] = 6'b000000;
		color_arr[1019] = 6'b000000;
		color_arr[1020] = 6'b000000;
		color_arr[1021] = 6'b000000;
		color_arr[1022] = 6'b000000;
		color_arr[1023] = 6'b000000;
		color_arr[1024] = 6'b000000;
		color_arr[1025] = 6'b000000;
		color_arr[1026] = 6'b000000;
		color_arr[1027] = 6'b000000;
		color_arr[1028] = 6'b000000;
		color_arr[1029] = 6'b000000;
		color_arr[1030] = 6'b000000;
		color_arr[1031] = 6'b000000;
		color_arr[1032] = 6'b000000;
		color_arr[1033] = 6'b000000;
		color_arr[1034] = 6'b000000;
		color_arr[1035] = 6'b000000;
		color_arr[1036] = 6'b000000;
		color_arr[1037] = 6'b000000;
		color_arr[1038] = 6'b000000;
		color_arr[1039] = 6'b000000;
		color_arr[1040] = 6'b111001;
		color_arr[1041] = 6'b111010;
		color_arr[1042] = 6'b111010;
		color_arr[1043] = 6'b111110;
		color_arr[1044] = 6'b111111;
		color_arr[1045] = 6'b000000;
		color_arr[1046] = 6'b000000;
		color_arr[1047] = 6'b111110;
		color_arr[1048] = 6'b111001;
		color_arr[1049] = 6'b111001;
		color_arr[1050] = 6'b111001;
		color_arr[1051] = 6'b111001;
		color_arr[1052] = 6'b111010;
		color_arr[1053] = 6'b111110;
		color_arr[1054] = 6'b111111;
		color_arr[1055] = 6'b111111;
		color_arr[1056] = 6'b111111;
		color_arr[1057] = 6'b111010;
		color_arr[1058] = 6'b111010;
		color_arr[1059] = 6'b111010;
		color_arr[1060] = 6'b111010;
		color_arr[1061] = 6'b111010;
		color_arr[1062] = 6'b111001;
		color_arr[1063] = 6'b111001;
		color_arr[1064] = 6'b111001;
		color_arr[1065] = 6'b000000;
		color_arr[1066] = 6'b000000;
		color_arr[1067] = 6'b000000;
		color_arr[1068] = 6'b000000;
		color_arr[1069] = 6'b000000;
		color_arr[1070] = 6'b000000;
		color_arr[1071] = 6'b000000;
		color_arr[1072] = 6'b000000;
		color_arr[1073] = 6'b000000;
		color_arr[1074] = 6'b000000;
		color_arr[1075] = 6'b000000;
		color_arr[1076] = 6'b000000;
		color_arr[1077] = 6'b000000;
		color_arr[1078] = 6'b000000;
		color_arr[1079] = 6'b000000;
		color_arr[1080] = 6'b000000;
		color_arr[1081] = 6'b000000;
		color_arr[1082] = 6'b000000;
		color_arr[1083] = 6'b000000;
		color_arr[1084] = 6'b000000;
		color_arr[1085] = 6'b000000;
		color_arr[1086] = 6'b000000;
		color_arr[1087] = 6'b000000;
		color_arr[1088] = 6'b000000;
		color_arr[1089] = 6'b000000;
		color_arr[1090] = 6'b000000;
		color_arr[1091] = 6'b000000;
		color_arr[1092] = 6'b000000;
		color_arr[1093] = 6'b000000;
		color_arr[1094] = 6'b000000;
		color_arr[1095] = 6'b000000;
		color_arr[1096] = 6'b000000;
		color_arr[1097] = 6'b000000;
		color_arr[1098] = 6'b000000;
		color_arr[1099] = 6'b000000;
		color_arr[1100] = 6'b000000;
		color_arr[1101] = 6'b000000;
		color_arr[1102] = 6'b000000;
		color_arr[1103] = 6'b000000;
		color_arr[1104] = 6'b111010;
		color_arr[1105] = 6'b111110;
		color_arr[1106] = 6'b111110;
		color_arr[1107] = 6'b111110;
		color_arr[1108] = 6'b111111;
		color_arr[1109] = 6'b000000;
		color_arr[1110] = 6'b000000;
		color_arr[1111] = 6'b111001;
		color_arr[1112] = 6'b111001;
		color_arr[1113] = 6'b111001;
		color_arr[1114] = 6'b111001;
		color_arr[1115] = 6'b111001;
		color_arr[1116] = 6'b111010;
		color_arr[1117] = 6'b111110;
		color_arr[1118] = 6'b111111;
		color_arr[1119] = 6'b000000;
		color_arr[1120] = 6'b000000;
		color_arr[1121] = 6'b111110;
		color_arr[1122] = 6'b111010;
		color_arr[1123] = 6'b111010;
		color_arr[1124] = 6'b111010;
		color_arr[1125] = 6'b111010;
		color_arr[1126] = 6'b111010;
		color_arr[1127] = 6'b111010;
		color_arr[1128] = 6'b111001;
		color_arr[1129] = 6'b111001;
		color_arr[1130] = 6'b000000;
		color_arr[1131] = 6'b000000;
		color_arr[1132] = 6'b000000;
		color_arr[1133] = 6'b000000;
		color_arr[1134] = 6'b000000;
		color_arr[1135] = 6'b000000;
		color_arr[1136] = 6'b000000;
		color_arr[1137] = 6'b000000;
		color_arr[1138] = 6'b000000;
		color_arr[1139] = 6'b000000;
		color_arr[1140] = 6'b000000;
		color_arr[1141] = 6'b000000;
		color_arr[1142] = 6'b000000;
		color_arr[1143] = 6'b000000;
		color_arr[1144] = 6'b000000;
		color_arr[1145] = 6'b000000;
		color_arr[1146] = 6'b000000;
		color_arr[1147] = 6'b000000;
		color_arr[1148] = 6'b000000;
		color_arr[1149] = 6'b000000;
		color_arr[1150] = 6'b000000;
		color_arr[1151] = 6'b000000;
		color_arr[1152] = 6'b000000;
		color_arr[1153] = 6'b000000;
		color_arr[1154] = 6'b000000;
		color_arr[1155] = 6'b000000;
		color_arr[1156] = 6'b000000;
		color_arr[1157] = 6'b000000;
		color_arr[1158] = 6'b000000;
		color_arr[1159] = 6'b000000;
		color_arr[1160] = 6'b000000;
		color_arr[1161] = 6'b000000;
		color_arr[1162] = 6'b000000;
		color_arr[1163] = 6'b000000;
		color_arr[1164] = 6'b000000;
		color_arr[1165] = 6'b000000;
		color_arr[1166] = 6'b000000;
		color_arr[1167] = 6'b111110;
		color_arr[1168] = 6'b111110;
		color_arr[1169] = 6'b111110;
		color_arr[1170] = 6'b111110;
		color_arr[1171] = 6'b111110;
		color_arr[1172] = 6'b111110;
		color_arr[1173] = 6'b111110;
		color_arr[1174] = 6'b111001;
		color_arr[1175] = 6'b111001;
		color_arr[1176] = 6'b111001;
		color_arr[1177] = 6'b111001;
		color_arr[1178] = 6'b111001;
		color_arr[1179] = 6'b111001;
		color_arr[1180] = 6'b111010;
		color_arr[1181] = 6'b111010;
		color_arr[1182] = 6'b111111;
		color_arr[1183] = 6'b000000;
		color_arr[1184] = 6'b000000;
		color_arr[1185] = 6'b111110;
		color_arr[1186] = 6'b111110;
		color_arr[1187] = 6'b111110;
		color_arr[1188] = 6'b111110;
		color_arr[1189] = 6'b111110;
		color_arr[1190] = 6'b111010;
		color_arr[1191] = 6'b111010;
		color_arr[1192] = 6'b111001;
		color_arr[1193] = 6'b111001;
		color_arr[1194] = 6'b000000;
		color_arr[1195] = 6'b000000;
		color_arr[1196] = 6'b000000;
		color_arr[1197] = 6'b000000;
		color_arr[1198] = 6'b000000;
		color_arr[1199] = 6'b000000;
		color_arr[1200] = 6'b000000;
		color_arr[1201] = 6'b000000;
		color_arr[1202] = 6'b000000;
		color_arr[1203] = 6'b000000;
		color_arr[1204] = 6'b000000;
		color_arr[1205] = 6'b000000;
		color_arr[1206] = 6'b000000;
		color_arr[1207] = 6'b000000;
		color_arr[1208] = 6'b000000;
		color_arr[1209] = 6'b000000;
		color_arr[1210] = 6'b000000;
		color_arr[1211] = 6'b000000;
		color_arr[1212] = 6'b000000;
		color_arr[1213] = 6'b000000;
		color_arr[1214] = 6'b000000;
		color_arr[1215] = 6'b000000;
		color_arr[1216] = 6'b000000;
		color_arr[1217] = 6'b000000;
		color_arr[1218] = 6'b000000;
		color_arr[1219] = 6'b000000;
		color_arr[1220] = 6'b000000;
		color_arr[1221] = 6'b000000;
		color_arr[1222] = 6'b000000;
		color_arr[1223] = 6'b000000;
		color_arr[1224] = 6'b000000;
		color_arr[1225] = 6'b000000;
		color_arr[1226] = 6'b000000;
		color_arr[1227] = 6'b000000;
		color_arr[1228] = 6'b000000;
		color_arr[1229] = 6'b000000;
		color_arr[1230] = 6'b000000;
		color_arr[1231] = 6'b111110;
		color_arr[1232] = 6'b111110;
		color_arr[1233] = 6'b111110;
		color_arr[1234] = 6'b111110;
		color_arr[1235] = 6'b111110;
		color_arr[1236] = 6'b111110;
		color_arr[1237] = 6'b111001;
		color_arr[1238] = 6'b111001;
		color_arr[1239] = 6'b111001;
		color_arr[1240] = 6'b111001;
		color_arr[1241] = 6'b111001;
		color_arr[1242] = 6'b111001;
		color_arr[1243] = 6'b111001;
		color_arr[1244] = 6'b111010;
		color_arr[1245] = 6'b111010;
		color_arr[1246] = 6'b111110;
		color_arr[1247] = 6'b111110;
		color_arr[1248] = 6'b111110;
		color_arr[1249] = 6'b111110;
		color_arr[1250] = 6'b111110;
		color_arr[1251] = 6'b111110;
		color_arr[1252] = 6'b111110;
		color_arr[1253] = 6'b111110;
		color_arr[1254] = 6'b111110;
		color_arr[1255] = 6'b111110;
		color_arr[1256] = 6'b111001;
		color_arr[1257] = 6'b111001;
		color_arr[1258] = 6'b111001;
		color_arr[1259] = 6'b000000;
		color_arr[1260] = 6'b000000;
		color_arr[1261] = 6'b000000;
		color_arr[1262] = 6'b000000;
		color_arr[1263] = 6'b000000;
		color_arr[1264] = 6'b000000;
		color_arr[1265] = 6'b000000;
		color_arr[1266] = 6'b000000;
		color_arr[1267] = 6'b000000;
		color_arr[1268] = 6'b000000;
		color_arr[1269] = 6'b000000;
		color_arr[1270] = 6'b000000;
		color_arr[1271] = 6'b000000;
		color_arr[1272] = 6'b000000;
		color_arr[1273] = 6'b000000;
		color_arr[1274] = 6'b000000;
		color_arr[1275] = 6'b000000;
		color_arr[1276] = 6'b000000;
		color_arr[1277] = 6'b000000;
		color_arr[1278] = 6'b000000;
		color_arr[1279] = 6'b000000;
		color_arr[1280] = 6'b000000;
		color_arr[1281] = 6'b000000;
		color_arr[1282] = 6'b000000;
		color_arr[1283] = 6'b000000;
		color_arr[1284] = 6'b000000;
		color_arr[1285] = 6'b000000;
		color_arr[1286] = 6'b000000;
		color_arr[1287] = 6'b000000;
		color_arr[1288] = 6'b000000;
		color_arr[1289] = 6'b000000;
		color_arr[1290] = 6'b000000;
		color_arr[1291] = 6'b000000;
		color_arr[1292] = 6'b000000;
		color_arr[1293] = 6'b000000;
		color_arr[1294] = 6'b000000;
		color_arr[1295] = 6'b111110;
		color_arr[1296] = 6'b111110;
		color_arr[1297] = 6'b111110;
		color_arr[1298] = 6'b111110;
		color_arr[1299] = 6'b111110;
		color_arr[1300] = 6'b111001;
		color_arr[1301] = 6'b111001;
		color_arr[1302] = 6'b111001;
		color_arr[1303] = 6'b111001;
		color_arr[1304] = 6'b111001;
		color_arr[1305] = 6'b111001;
		color_arr[1306] = 6'b111001;
		color_arr[1307] = 6'b111001;
		color_arr[1308] = 6'b111010;
		color_arr[1309] = 6'b111010;
		color_arr[1310] = 6'b111010;
		color_arr[1311] = 6'b111110;
		color_arr[1312] = 6'b111110;
		color_arr[1313] = 6'b111110;
		color_arr[1314] = 6'b111110;
		color_arr[1315] = 6'b111110;
		color_arr[1316] = 6'b111110;
		color_arr[1317] = 6'b111110;
		color_arr[1318] = 6'b111110;
		color_arr[1319] = 6'b111110;
		color_arr[1320] = 6'b111110;
		color_arr[1321] = 6'b111001;
		color_arr[1322] = 6'b111001;
		color_arr[1323] = 6'b000000;
		color_arr[1324] = 6'b000000;
		color_arr[1325] = 6'b000000;
		color_arr[1326] = 6'b000000;
		color_arr[1327] = 6'b000000;
		color_arr[1328] = 6'b000000;
		color_arr[1329] = 6'b000000;
		color_arr[1330] = 6'b000000;
		color_arr[1331] = 6'b000000;
		color_arr[1332] = 6'b000000;
		color_arr[1333] = 6'b000000;
		color_arr[1334] = 6'b000000;
		color_arr[1335] = 6'b000000;
		color_arr[1336] = 6'b000000;
		color_arr[1337] = 6'b000000;
		color_arr[1338] = 6'b000000;
		color_arr[1339] = 6'b000000;
		color_arr[1340] = 6'b000000;
		color_arr[1341] = 6'b000000;
		color_arr[1342] = 6'b000000;
		color_arr[1343] = 6'b000000;
		color_arr[1344] = 6'b000000;
		color_arr[1345] = 6'b000000;
		color_arr[1346] = 6'b000000;
		color_arr[1347] = 6'b000000;
		color_arr[1348] = 6'b000000;
		color_arr[1349] = 6'b000000;
		color_arr[1350] = 6'b000000;
		color_arr[1351] = 6'b000000;
		color_arr[1352] = 6'b000000;
		color_arr[1353] = 6'b000000;
		color_arr[1354] = 6'b000000;
		color_arr[1355] = 6'b000000;
		color_arr[1356] = 6'b000000;
		color_arr[1357] = 6'b000000;
		color_arr[1358] = 6'b000000;
		color_arr[1359] = 6'b111110;
		color_arr[1360] = 6'b111110;
		color_arr[1361] = 6'b111110;
		color_arr[1362] = 6'b111110;
		color_arr[1363] = 6'b010101;
		color_arr[1364] = 6'b010101;
		color_arr[1365] = 6'b000000;
		color_arr[1366] = 6'b000000;
		color_arr[1367] = 6'b000000;
		color_arr[1368] = 6'b111111;
		color_arr[1369] = 6'b111001;
		color_arr[1370] = 6'b111001;
		color_arr[1371] = 6'b111010;
		color_arr[1372] = 6'b111010;
		color_arr[1373] = 6'b111010;
		color_arr[1374] = 6'b111110;
		color_arr[1375] = 6'b111110;
		color_arr[1376] = 6'b111110;
		color_arr[1377] = 6'b111110;
		color_arr[1378] = 6'b111110;
		color_arr[1379] = 6'b111110;
		color_arr[1380] = 6'b111110;
		color_arr[1381] = 6'b111110;
		color_arr[1382] = 6'b111110;
		color_arr[1383] = 6'b111110;
		color_arr[1384] = 6'b111110;
		color_arr[1385] = 6'b111001;
		color_arr[1386] = 6'b111001;
		color_arr[1387] = 6'b111001;
		color_arr[1388] = 6'b000000;
		color_arr[1389] = 6'b000000;
		color_arr[1390] = 6'b000000;
		color_arr[1391] = 6'b000000;
		color_arr[1392] = 6'b000000;
		color_arr[1393] = 6'b000000;
		color_arr[1394] = 6'b000000;
		color_arr[1395] = 6'b000000;
		color_arr[1396] = 6'b000000;
		color_arr[1397] = 6'b000000;
		color_arr[1398] = 6'b000000;
		color_arr[1399] = 6'b000000;
		color_arr[1400] = 6'b000000;
		color_arr[1401] = 6'b000000;
		color_arr[1402] = 6'b000000;
		color_arr[1403] = 6'b000000;
		color_arr[1404] = 6'b000000;
		color_arr[1405] = 6'b000000;
		color_arr[1406] = 6'b000000;
		color_arr[1407] = 6'b000000;
		color_arr[1408] = 6'b000000;
		color_arr[1409] = 6'b000000;
		color_arr[1410] = 6'b000000;
		color_arr[1411] = 6'b000000;
		color_arr[1412] = 6'b000000;
		color_arr[1413] = 6'b000000;
		color_arr[1414] = 6'b000000;
		color_arr[1415] = 6'b000000;
		color_arr[1416] = 6'b000000;
		color_arr[1417] = 6'b000000;
		color_arr[1418] = 6'b000000;
		color_arr[1419] = 6'b000000;
		color_arr[1420] = 6'b000000;
		color_arr[1421] = 6'b000000;
		color_arr[1422] = 6'b000000;
		color_arr[1423] = 6'b111110;
		color_arr[1424] = 6'b111110;
		color_arr[1425] = 6'b111110;
		color_arr[1426] = 6'b111110;
		color_arr[1427] = 6'b010101;
		color_arr[1428] = 6'b000000;
		color_arr[1429] = 6'b000000;
		color_arr[1430] = 6'b000000;
		color_arr[1431] = 6'b000000;
		color_arr[1432] = 6'b111111;
		color_arr[1433] = 6'b111111;
		color_arr[1434] = 6'b111010;
		color_arr[1435] = 6'b111010;
		color_arr[1436] = 6'b111010;
		color_arr[1437] = 6'b111010;
		color_arr[1438] = 6'b111110;
		color_arr[1439] = 6'b111110;
		color_arr[1440] = 6'b111110;
		color_arr[1441] = 6'b111110;
		color_arr[1442] = 6'b111110;
		color_arr[1443] = 6'b111110;
		color_arr[1444] = 6'b111110;
		color_arr[1445] = 6'b111110;
		color_arr[1446] = 6'b111110;
		color_arr[1447] = 6'b111110;
		color_arr[1448] = 6'b111110;
		color_arr[1449] = 6'b111001;
		color_arr[1450] = 6'b111001;
		color_arr[1451] = 6'b111001;
		color_arr[1452] = 6'b000000;
		color_arr[1453] = 6'b000000;
		color_arr[1454] = 6'b000000;
		color_arr[1455] = 6'b000000;
		color_arr[1456] = 6'b000000;
		color_arr[1457] = 6'b000000;
		color_arr[1458] = 6'b000000;
		color_arr[1459] = 6'b000000;
		color_arr[1460] = 6'b000000;
		color_arr[1461] = 6'b000000;
		color_arr[1462] = 6'b000000;
		color_arr[1463] = 6'b000000;
		color_arr[1464] = 6'b000000;
		color_arr[1465] = 6'b000000;
		color_arr[1466] = 6'b000000;
		color_arr[1467] = 6'b000000;
		color_arr[1468] = 6'b000000;
		color_arr[1469] = 6'b000000;
		color_arr[1470] = 6'b000000;
		color_arr[1471] = 6'b000000;
		color_arr[1472] = 6'b000000;
		color_arr[1473] = 6'b000000;
		color_arr[1474] = 6'b000000;
		color_arr[1475] = 6'b000000;
		color_arr[1476] = 6'b000000;
		color_arr[1477] = 6'b000000;
		color_arr[1478] = 6'b000000;
		color_arr[1479] = 6'b000000;
		color_arr[1480] = 6'b000000;
		color_arr[1481] = 6'b000000;
		color_arr[1482] = 6'b000000;
		color_arr[1483] = 6'b000000;
		color_arr[1484] = 6'b000000;
		color_arr[1485] = 6'b000000;
		color_arr[1486] = 6'b000000;
		color_arr[1487] = 6'b111110;
		color_arr[1488] = 6'b111110;
		color_arr[1489] = 6'b111110;
		color_arr[1490] = 6'b111111;
		color_arr[1491] = 6'b111111;
		color_arr[1492] = 6'b000000;
		color_arr[1493] = 6'b000000;
		color_arr[1494] = 6'b000000;
		color_arr[1495] = 6'b111111;
		color_arr[1496] = 6'b111111;
		color_arr[1497] = 6'b111111;
		color_arr[1498] = 6'b111111;
		color_arr[1499] = 6'b111111;
		color_arr[1500] = 6'b111010;
		color_arr[1501] = 6'b111110;
		color_arr[1502] = 6'b111110;
		color_arr[1503] = 6'b111110;
		color_arr[1504] = 6'b111110;
		color_arr[1505] = 6'b111110;
		color_arr[1506] = 6'b111110;
		color_arr[1507] = 6'b111110;
		color_arr[1508] = 6'b111110;
		color_arr[1509] = 6'b111110;
		color_arr[1510] = 6'b111110;
		color_arr[1511] = 6'b111110;
		color_arr[1512] = 6'b111110;
		color_arr[1513] = 6'b111110;
		color_arr[1514] = 6'b111001;
		color_arr[1515] = 6'b111001;
		color_arr[1516] = 6'b000000;
		color_arr[1517] = 6'b000000;
		color_arr[1518] = 6'b000000;
		color_arr[1519] = 6'b000000;
		color_arr[1520] = 6'b000000;
		color_arr[1521] = 6'b000000;
		color_arr[1522] = 6'b000000;
		color_arr[1523] = 6'b000000;
		color_arr[1524] = 6'b000000;
		color_arr[1525] = 6'b000000;
		color_arr[1526] = 6'b000000;
		color_arr[1527] = 6'b000000;
		color_arr[1528] = 6'b000000;
		color_arr[1529] = 6'b000000;
		color_arr[1530] = 6'b000000;
		color_arr[1531] = 6'b000000;
		color_arr[1532] = 6'b000000;
		color_arr[1533] = 6'b000000;
		color_arr[1534] = 6'b000000;
		color_arr[1535] = 6'b000000;
		color_arr[1536] = 6'b000000;
		color_arr[1537] = 6'b000000;
		color_arr[1538] = 6'b000000;
		color_arr[1539] = 6'b000000;
		color_arr[1540] = 6'b000000;
		color_arr[1541] = 6'b000000;
		color_arr[1542] = 6'b000000;
		color_arr[1543] = 6'b000000;
		color_arr[1544] = 6'b000000;
		color_arr[1545] = 6'b000000;
		color_arr[1546] = 6'b000000;
		color_arr[1547] = 6'b000000;
		color_arr[1548] = 6'b000000;
		color_arr[1549] = 6'b000000;
		color_arr[1550] = 6'b000000;
		color_arr[1551] = 6'b111110;
		color_arr[1552] = 6'b111110;
		color_arr[1553] = 6'b111110;
		color_arr[1554] = 6'b111111;
		color_arr[1555] = 6'b010101;
		color_arr[1556] = 6'b010101;
		color_arr[1557] = 6'b000000;
		color_arr[1558] = 6'b010101;
		color_arr[1559] = 6'b111111;
		color_arr[1560] = 6'b111111;
		color_arr[1561] = 6'b111111;
		color_arr[1562] = 6'b111111;
		color_arr[1563] = 6'b111111;
		color_arr[1564] = 6'b111111;
		color_arr[1565] = 6'b000000;
		color_arr[1566] = 6'b111110;
		color_arr[1567] = 6'b111110;
		color_arr[1568] = 6'b111110;
		color_arr[1569] = 6'b111110;
		color_arr[1570] = 6'b111110;
		color_arr[1571] = 6'b111110;
		color_arr[1572] = 6'b111110;
		color_arr[1573] = 6'b111110;
		color_arr[1574] = 6'b111110;
		color_arr[1575] = 6'b111110;
		color_arr[1576] = 6'b111110;
		color_arr[1577] = 6'b111110;
		color_arr[1578] = 6'b111001;
		color_arr[1579] = 6'b111001;
		color_arr[1580] = 6'b000000;
		color_arr[1581] = 6'b000000;
		color_arr[1582] = 6'b000000;
		color_arr[1583] = 6'b000000;
		color_arr[1584] = 6'b000000;
		color_arr[1585] = 6'b000000;
		color_arr[1586] = 6'b000000;
		color_arr[1587] = 6'b000000;
		color_arr[1588] = 6'b000000;
		color_arr[1589] = 6'b000000;
		color_arr[1590] = 6'b000000;
		color_arr[1591] = 6'b000000;
		color_arr[1592] = 6'b000000;
		color_arr[1593] = 6'b000000;
		color_arr[1594] = 6'b000000;
		color_arr[1595] = 6'b000000;
		color_arr[1596] = 6'b000000;
		color_arr[1597] = 6'b000000;
		color_arr[1598] = 6'b000000;
		color_arr[1599] = 6'b000000;
		color_arr[1600] = 6'b000000;
		color_arr[1601] = 6'b000000;
		color_arr[1602] = 6'b000000;
		color_arr[1603] = 6'b000000;
		color_arr[1604] = 6'b000000;
		color_arr[1605] = 6'b000000;
		color_arr[1606] = 6'b000000;
		color_arr[1607] = 6'b000000;
		color_arr[1608] = 6'b000000;
		color_arr[1609] = 6'b000000;
		color_arr[1610] = 6'b000000;
		color_arr[1611] = 6'b000000;
		color_arr[1612] = 6'b000000;
		color_arr[1613] = 6'b000000;
		color_arr[1614] = 6'b000000;
		color_arr[1615] = 6'b000000;
		color_arr[1616] = 6'b111110;
		color_arr[1617] = 6'b111110;
		color_arr[1618] = 6'b111110;
		color_arr[1619] = 6'b000000;
		color_arr[1620] = 6'b000000;
		color_arr[1621] = 6'b010101;
		color_arr[1622] = 6'b010101;
		color_arr[1623] = 6'b010101;
		color_arr[1624] = 6'b010101;
		color_arr[1625] = 6'b111111;
		color_arr[1626] = 6'b111111;
		color_arr[1627] = 6'b000000;
		color_arr[1628] = 6'b000000;
		color_arr[1629] = 6'b111110;
		color_arr[1630] = 6'b111110;
		color_arr[1631] = 6'b111110;
		color_arr[1632] = 6'b111110;
		color_arr[1633] = 6'b111110;
		color_arr[1634] = 6'b111110;
		color_arr[1635] = 6'b111110;
		color_arr[1636] = 6'b111110;
		color_arr[1637] = 6'b111110;
		color_arr[1638] = 6'b111110;
		color_arr[1639] = 6'b111110;
		color_arr[1640] = 6'b111110;
		color_arr[1641] = 6'b111110;
		color_arr[1642] = 6'b111001;
		color_arr[1643] = 6'b111001;
		color_arr[1644] = 6'b111001;
		color_arr[1645] = 6'b000000;
		color_arr[1646] = 6'b000000;
		color_arr[1647] = 6'b000000;
		color_arr[1648] = 6'b000000;
		color_arr[1649] = 6'b000000;
		color_arr[1650] = 6'b000000;
		color_arr[1651] = 6'b000000;
		color_arr[1652] = 6'b000000;
		color_arr[1653] = 6'b000000;
		color_arr[1654] = 6'b000000;
		color_arr[1655] = 6'b000000;
		color_arr[1656] = 6'b000000;
		color_arr[1657] = 6'b000000;
		color_arr[1658] = 6'b000000;
		color_arr[1659] = 6'b000000;
		color_arr[1660] = 6'b000000;
		color_arr[1661] = 6'b000000;
		color_arr[1662] = 6'b000000;
		color_arr[1663] = 6'b000000;
		color_arr[1664] = 6'b000000;
		color_arr[1665] = 6'b000000;
		color_arr[1666] = 6'b000000;
		color_arr[1667] = 6'b000000;
		color_arr[1668] = 6'b000000;
		color_arr[1669] = 6'b000000;
		color_arr[1670] = 6'b000000;
		color_arr[1671] = 6'b000000;
		color_arr[1672] = 6'b000000;
		color_arr[1673] = 6'b000000;
		color_arr[1674] = 6'b000000;
		color_arr[1675] = 6'b000000;
		color_arr[1676] = 6'b000000;
		color_arr[1677] = 6'b000000;
		color_arr[1678] = 6'b000000;
		color_arr[1679] = 6'b000000;
		color_arr[1680] = 6'b111110;
		color_arr[1681] = 6'b111110;
		color_arr[1682] = 6'b111110;
		color_arr[1683] = 6'b111110;
		color_arr[1684] = 6'b111110;
		color_arr[1685] = 6'b000000;
		color_arr[1686] = 6'b000000;
		color_arr[1687] = 6'b000000;
		color_arr[1688] = 6'b000000;
		color_arr[1689] = 6'b000000;
		color_arr[1690] = 6'b000000;
		color_arr[1691] = 6'b111110;
		color_arr[1692] = 6'b111110;
		color_arr[1693] = 6'b111110;
		color_arr[1694] = 6'b111110;
		color_arr[1695] = 6'b111110;
		color_arr[1696] = 6'b111110;
		color_arr[1697] = 6'b111110;
		color_arr[1698] = 6'b111110;
		color_arr[1699] = 6'b111110;
		color_arr[1700] = 6'b111110;
		color_arr[1701] = 6'b111110;
		color_arr[1702] = 6'b111110;
		color_arr[1703] = 6'b111110;
		color_arr[1704] = 6'b111110;
		color_arr[1705] = 6'b111110;
		color_arr[1706] = 6'b111010;
		color_arr[1707] = 6'b111001;
		color_arr[1708] = 6'b111001;
		color_arr[1709] = 6'b000000;
		color_arr[1710] = 6'b000000;
		color_arr[1711] = 6'b000000;
		color_arr[1712] = 6'b000000;
		color_arr[1713] = 6'b000000;
		color_arr[1714] = 6'b000000;
		color_arr[1715] = 6'b000000;
		color_arr[1716] = 6'b000000;
		color_arr[1717] = 6'b000000;
		color_arr[1718] = 6'b000000;
		color_arr[1719] = 6'b000000;
		color_arr[1720] = 6'b000000;
		color_arr[1721] = 6'b000000;
		color_arr[1722] = 6'b000000;
		color_arr[1723] = 6'b000000;
		color_arr[1724] = 6'b000000;
		color_arr[1725] = 6'b000000;
		color_arr[1726] = 6'b000000;
		color_arr[1727] = 6'b000000;
		color_arr[1728] = 6'b000000;
		color_arr[1729] = 6'b000000;
		color_arr[1730] = 6'b000000;
		color_arr[1731] = 6'b000000;
		color_arr[1732] = 6'b000000;
		color_arr[1733] = 6'b000000;
		color_arr[1734] = 6'b000000;
		color_arr[1735] = 6'b000000;
		color_arr[1736] = 6'b000000;
		color_arr[1737] = 6'b000000;
		color_arr[1738] = 6'b000000;
		color_arr[1739] = 6'b000000;
		color_arr[1740] = 6'b000000;
		color_arr[1741] = 6'b000000;
		color_arr[1742] = 6'b000000;
		color_arr[1743] = 6'b000000;
		color_arr[1744] = 6'b000000;
		color_arr[1745] = 6'b111110;
		color_arr[1746] = 6'b111110;
		color_arr[1747] = 6'b111110;
		color_arr[1748] = 6'b111110;
		color_arr[1749] = 6'b111110;
		color_arr[1750] = 6'b111110;
		color_arr[1751] = 6'b111110;
		color_arr[1752] = 6'b111110;
		color_arr[1753] = 6'b111110;
		color_arr[1754] = 6'b111110;
		color_arr[1755] = 6'b111110;
		color_arr[1756] = 6'b111110;
		color_arr[1757] = 6'b111110;
		color_arr[1758] = 6'b111110;
		color_arr[1759] = 6'b111110;
		color_arr[1760] = 6'b111110;
		color_arr[1761] = 6'b111110;
		color_arr[1762] = 6'b111110;
		color_arr[1763] = 6'b111110;
		color_arr[1764] = 6'b111110;
		color_arr[1765] = 6'b111110;
		color_arr[1766] = 6'b111110;
		color_arr[1767] = 6'b111110;
		color_arr[1768] = 6'b111110;
		color_arr[1769] = 6'b111110;
		color_arr[1770] = 6'b111010;
		color_arr[1771] = 6'b111001;
		color_arr[1772] = 6'b111001;
		color_arr[1773] = 6'b000000;
		color_arr[1774] = 6'b000000;
		color_arr[1775] = 6'b000000;
		color_arr[1776] = 6'b000000;
		color_arr[1777] = 6'b000000;
		color_arr[1778] = 6'b000000;
		color_arr[1779] = 6'b000000;
		color_arr[1780] = 6'b000000;
		color_arr[1781] = 6'b000000;
		color_arr[1782] = 6'b000000;
		color_arr[1783] = 6'b000000;
		color_arr[1784] = 6'b000000;
		color_arr[1785] = 6'b000000;
		color_arr[1786] = 6'b000000;
		color_arr[1787] = 6'b000000;
		color_arr[1788] = 6'b000000;
		color_arr[1789] = 6'b000000;
		color_arr[1790] = 6'b000000;
		color_arr[1791] = 6'b000000;
		color_arr[1792] = 6'b000000;
		color_arr[1793] = 6'b000000;
		color_arr[1794] = 6'b000000;
		color_arr[1795] = 6'b000000;
		color_arr[1796] = 6'b000000;
		color_arr[1797] = 6'b000000;
		color_arr[1798] = 6'b000000;
		color_arr[1799] = 6'b000000;
		color_arr[1800] = 6'b000000;
		color_arr[1801] = 6'b000000;
		color_arr[1802] = 6'b000000;
		color_arr[1803] = 6'b000000;
		color_arr[1804] = 6'b000000;
		color_arr[1805] = 6'b000000;
		color_arr[1806] = 6'b000000;
		color_arr[1807] = 6'b000000;
		color_arr[1808] = 6'b000000;
		color_arr[1809] = 6'b000000;
		color_arr[1810] = 6'b111110;
		color_arr[1811] = 6'b111110;
		color_arr[1812] = 6'b111110;
		color_arr[1813] = 6'b111110;
		color_arr[1814] = 6'b111110;
		color_arr[1815] = 6'b111110;
		color_arr[1816] = 6'b111110;
		color_arr[1817] = 6'b111110;
		color_arr[1818] = 6'b111110;
		color_arr[1819] = 6'b111110;
		color_arr[1820] = 6'b111110;
		color_arr[1821] = 6'b111110;
		color_arr[1822] = 6'b111110;
		color_arr[1823] = 6'b111110;
		color_arr[1824] = 6'b111110;
		color_arr[1825] = 6'b111110;
		color_arr[1826] = 6'b111110;
		color_arr[1827] = 6'b111110;
		color_arr[1828] = 6'b111110;
		color_arr[1829] = 6'b111110;
		color_arr[1830] = 6'b111110;
		color_arr[1831] = 6'b111110;
		color_arr[1832] = 6'b111110;
		color_arr[1833] = 6'b111010;
		color_arr[1834] = 6'b111010;
		color_arr[1835] = 6'b111010;
		color_arr[1836] = 6'b111001;
		color_arr[1837] = 6'b111001;
		color_arr[1838] = 6'b000000;
		color_arr[1839] = 6'b000000;
		color_arr[1840] = 6'b000000;
		color_arr[1841] = 6'b000000;
		color_arr[1842] = 6'b000000;
		color_arr[1843] = 6'b000000;
		color_arr[1844] = 6'b000000;
		color_arr[1845] = 6'b000000;
		color_arr[1846] = 6'b000000;
		color_arr[1847] = 6'b000000;
		color_arr[1848] = 6'b000000;
		color_arr[1849] = 6'b000000;
		color_arr[1850] = 6'b000000;
		color_arr[1851] = 6'b000000;
		color_arr[1852] = 6'b000000;
		color_arr[1853] = 6'b000000;
		color_arr[1854] = 6'b000000;
		color_arr[1855] = 6'b000000;
		color_arr[1856] = 6'b000000;
		color_arr[1857] = 6'b000000;
		color_arr[1858] = 6'b000000;
		color_arr[1859] = 6'b000000;
		color_arr[1860] = 6'b000000;
		color_arr[1861] = 6'b000000;
		color_arr[1862] = 6'b000000;
		color_arr[1863] = 6'b000000;
		color_arr[1864] = 6'b000000;
		color_arr[1865] = 6'b000000;
		color_arr[1866] = 6'b000000;
		color_arr[1867] = 6'b000000;
		color_arr[1868] = 6'b000000;
		color_arr[1869] = 6'b000000;
		color_arr[1870] = 6'b000000;
		color_arr[1871] = 6'b000000;
		color_arr[1872] = 6'b000000;
		color_arr[1873] = 6'b000000;
		color_arr[1874] = 6'b111110;
		color_arr[1875] = 6'b111110;
		color_arr[1876] = 6'b111110;
		color_arr[1877] = 6'b111110;
		color_arr[1878] = 6'b111110;
		color_arr[1879] = 6'b111110;
		color_arr[1880] = 6'b111110;
		color_arr[1881] = 6'b111110;
		color_arr[1882] = 6'b111110;
		color_arr[1883] = 6'b111110;
		color_arr[1884] = 6'b111110;
		color_arr[1885] = 6'b111110;
		color_arr[1886] = 6'b111110;
		color_arr[1887] = 6'b111110;
		color_arr[1888] = 6'b111110;
		color_arr[1889] = 6'b111110;
		color_arr[1890] = 6'b111110;
		color_arr[1891] = 6'b111110;
		color_arr[1892] = 6'b111110;
		color_arr[1893] = 6'b111110;
		color_arr[1894] = 6'b111110;
		color_arr[1895] = 6'b111110;
		color_arr[1896] = 6'b111010;
		color_arr[1897] = 6'b111010;
		color_arr[1898] = 6'b111001;
		color_arr[1899] = 6'b111010;
		color_arr[1900] = 6'b111001;
		color_arr[1901] = 6'b111001;
		color_arr[1902] = 6'b000000;
		color_arr[1903] = 6'b000000;
		color_arr[1904] = 6'b000000;
		color_arr[1905] = 6'b000000;
		color_arr[1906] = 6'b000000;
		color_arr[1907] = 6'b000000;
		color_arr[1908] = 6'b000000;
		color_arr[1909] = 6'b000000;
		color_arr[1910] = 6'b000000;
		color_arr[1911] = 6'b000000;
		color_arr[1912] = 6'b000000;
		color_arr[1913] = 6'b000000;
		color_arr[1914] = 6'b000000;
		color_arr[1915] = 6'b000000;
		color_arr[1916] = 6'b000000;
		color_arr[1917] = 6'b000000;
		color_arr[1918] = 6'b000000;
		color_arr[1919] = 6'b000000;
		color_arr[1920] = 6'b000000;
		color_arr[1921] = 6'b000000;
		color_arr[1922] = 6'b000000;
		color_arr[1923] = 6'b000000;
		color_arr[1924] = 6'b000000;
		color_arr[1925] = 6'b000000;
		color_arr[1926] = 6'b000000;
		color_arr[1927] = 6'b000000;
		color_arr[1928] = 6'b000000;
		color_arr[1929] = 6'b000000;
		color_arr[1930] = 6'b000000;
		color_arr[1931] = 6'b000000;
		color_arr[1932] = 6'b000000;
		color_arr[1933] = 6'b000000;
		color_arr[1934] = 6'b000000;
		color_arr[1935] = 6'b000000;
		color_arr[1936] = 6'b000000;
		color_arr[1937] = 6'b000000;
		color_arr[1938] = 6'b000000;
		color_arr[1939] = 6'b111110;
		color_arr[1940] = 6'b111110;
		color_arr[1941] = 6'b111110;
		color_arr[1942] = 6'b111110;
		color_arr[1943] = 6'b111110;
		color_arr[1944] = 6'b111110;
		color_arr[1945] = 6'b111110;
		color_arr[1946] = 6'b111110;
		color_arr[1947] = 6'b111110;
		color_arr[1948] = 6'b111110;
		color_arr[1949] = 6'b111110;
		color_arr[1950] = 6'b111110;
		color_arr[1951] = 6'b111110;
		color_arr[1952] = 6'b111110;
		color_arr[1953] = 6'b111110;
		color_arr[1954] = 6'b111110;
		color_arr[1955] = 6'b111110;
		color_arr[1956] = 6'b111110;
		color_arr[1957] = 6'b111110;
		color_arr[1958] = 6'b111110;
		color_arr[1959] = 6'b111010;
		color_arr[1960] = 6'b111010;
		color_arr[1961] = 6'b111001;
		color_arr[1962] = 6'b111001;
		color_arr[1963] = 6'b111010;
		color_arr[1964] = 6'b111001;
		color_arr[1965] = 6'b111001;
		color_arr[1966] = 6'b111001;
		color_arr[1967] = 6'b000000;
		color_arr[1968] = 6'b000000;
		color_arr[1969] = 6'b000000;
		color_arr[1970] = 6'b000000;
		color_arr[1971] = 6'b000000;
		color_arr[1972] = 6'b000000;
		color_arr[1973] = 6'b000000;
		color_arr[1974] = 6'b000000;
		color_arr[1975] = 6'b000000;
		color_arr[1976] = 6'b000000;
		color_arr[1977] = 6'b000000;
		color_arr[1978] = 6'b000000;
		color_arr[1979] = 6'b000000;
		color_arr[1980] = 6'b000000;
		color_arr[1981] = 6'b000000;
		color_arr[1982] = 6'b000000;
		color_arr[1983] = 6'b000000;
		color_arr[1984] = 6'b000000;
		color_arr[1985] = 6'b000000;
		color_arr[1986] = 6'b000000;
		color_arr[1987] = 6'b000000;
		color_arr[1988] = 6'b000000;
		color_arr[1989] = 6'b000000;
		color_arr[1990] = 6'b000000;
		color_arr[1991] = 6'b000000;
		color_arr[1992] = 6'b000000;
		color_arr[1993] = 6'b000000;
		color_arr[1994] = 6'b000000;
		color_arr[1995] = 6'b000000;
		color_arr[1996] = 6'b000000;
		color_arr[1997] = 6'b000000;
		color_arr[1998] = 6'b000000;
		color_arr[1999] = 6'b000000;
		color_arr[2000] = 6'b000000;
		color_arr[2001] = 6'b000000;
		color_arr[2002] = 6'b000000;
		color_arr[2003] = 6'b111110;
		color_arr[2004] = 6'b111110;
		color_arr[2005] = 6'b111110;
		color_arr[2006] = 6'b111110;
		color_arr[2007] = 6'b111110;
		color_arr[2008] = 6'b111110;
		color_arr[2009] = 6'b111110;
		color_arr[2010] = 6'b111110;
		color_arr[2011] = 6'b111110;
		color_arr[2012] = 6'b111110;
		color_arr[2013] = 6'b111110;
		color_arr[2014] = 6'b111110;
		color_arr[2015] = 6'b111110;
		color_arr[2016] = 6'b111110;
		color_arr[2017] = 6'b111110;
		color_arr[2018] = 6'b111110;
		color_arr[2019] = 6'b111110;
		color_arr[2020] = 6'b111110;
		color_arr[2021] = 6'b111110;
		color_arr[2022] = 6'b111010;
		color_arr[2023] = 6'b111010;
		color_arr[2024] = 6'b111001;
		color_arr[2025] = 6'b111001;
		color_arr[2026] = 6'b111001;
		color_arr[2027] = 6'b111010;
		color_arr[2028] = 6'b111001;
		color_arr[2029] = 6'b111001;
		color_arr[2030] = 6'b111001;
		color_arr[2031] = 6'b000000;
		color_arr[2032] = 6'b000000;
		color_arr[2033] = 6'b000000;
		color_arr[2034] = 6'b000000;
		color_arr[2035] = 6'b000000;
		color_arr[2036] = 6'b000000;
		color_arr[2037] = 6'b000000;
		color_arr[2038] = 6'b000000;
		color_arr[2039] = 6'b000000;
		color_arr[2040] = 6'b000000;
		color_arr[2041] = 6'b000000;
		color_arr[2042] = 6'b000000;
		color_arr[2043] = 6'b000000;
		color_arr[2044] = 6'b000000;
		color_arr[2045] = 6'b000000;
		color_arr[2046] = 6'b000000;
		color_arr[2047] = 6'b000000;
		color_arr[2048] = 6'b000000;
		color_arr[2049] = 6'b000000;
		color_arr[2050] = 6'b000000;
		color_arr[2051] = 6'b000000;
		color_arr[2052] = 6'b000000;
		color_arr[2053] = 6'b000000;
		color_arr[2054] = 6'b000000;
		color_arr[2055] = 6'b000000;
		color_arr[2056] = 6'b000000;
		color_arr[2057] = 6'b000000;
		color_arr[2058] = 6'b000000;
		color_arr[2059] = 6'b000000;
		color_arr[2060] = 6'b000000;
		color_arr[2061] = 6'b000000;
		color_arr[2062] = 6'b000000;
		color_arr[2063] = 6'b000000;
		color_arr[2064] = 6'b000000;
		color_arr[2065] = 6'b000000;
		color_arr[2066] = 6'b000000;
		color_arr[2067] = 6'b000000;
		color_arr[2068] = 6'b111110;
		color_arr[2069] = 6'b111110;
		color_arr[2070] = 6'b111110;
		color_arr[2071] = 6'b111110;
		color_arr[2072] = 6'b111110;
		color_arr[2073] = 6'b111110;
		color_arr[2074] = 6'b111110;
		color_arr[2075] = 6'b111110;
		color_arr[2076] = 6'b111110;
		color_arr[2077] = 6'b111110;
		color_arr[2078] = 6'b111110;
		color_arr[2079] = 6'b111110;
		color_arr[2080] = 6'b111110;
		color_arr[2081] = 6'b111110;
		color_arr[2082] = 6'b111110;
		color_arr[2083] = 6'b111110;
		color_arr[2084] = 6'b111110;
		color_arr[2085] = 6'b111010;
		color_arr[2086] = 6'b111010;
		color_arr[2087] = 6'b111001;
		color_arr[2088] = 6'b111001;
		color_arr[2089] = 6'b111001;
		color_arr[2090] = 6'b111001;
		color_arr[2091] = 6'b111010;
		color_arr[2092] = 6'b111010;
		color_arr[2093] = 6'b111001;
		color_arr[2094] = 6'b111001;
		color_arr[2095] = 6'b000000;
		color_arr[2096] = 6'b000000;
		color_arr[2097] = 6'b000000;
		color_arr[2098] = 6'b000000;
		color_arr[2099] = 6'b000000;
		color_arr[2100] = 6'b000000;
		color_arr[2101] = 6'b000000;
		color_arr[2102] = 6'b000000;
		color_arr[2103] = 6'b000000;
		color_arr[2104] = 6'b000000;
		color_arr[2105] = 6'b000000;
		color_arr[2106] = 6'b000000;
		color_arr[2107] = 6'b000000;
		color_arr[2108] = 6'b000000;
		color_arr[2109] = 6'b000000;
		color_arr[2110] = 6'b000000;
		color_arr[2111] = 6'b000000;
		color_arr[2112] = 6'b000000;
		color_arr[2113] = 6'b000000;
		color_arr[2114] = 6'b000000;
		color_arr[2115] = 6'b000000;
		color_arr[2116] = 6'b000000;
		color_arr[2117] = 6'b000000;
		color_arr[2118] = 6'b000000;
		color_arr[2119] = 6'b000000;
		color_arr[2120] = 6'b000000;
		color_arr[2121] = 6'b000000;
		color_arr[2122] = 6'b000000;
		color_arr[2123] = 6'b000000;
		color_arr[2124] = 6'b000000;
		color_arr[2125] = 6'b000000;
		color_arr[2126] = 6'b000000;
		color_arr[2127] = 6'b000000;
		color_arr[2128] = 6'b000000;
		color_arr[2129] = 6'b000000;
		color_arr[2130] = 6'b000000;
		color_arr[2131] = 6'b000000;
		color_arr[2132] = 6'b111110;
		color_arr[2133] = 6'b111110;
		color_arr[2134] = 6'b111110;
		color_arr[2135] = 6'b111110;
		color_arr[2136] = 6'b111110;
		color_arr[2137] = 6'b111110;
		color_arr[2138] = 6'b111110;
		color_arr[2139] = 6'b111110;
		color_arr[2140] = 6'b111110;
		color_arr[2141] = 6'b111110;
		color_arr[2142] = 6'b111110;
		color_arr[2143] = 6'b111110;
		color_arr[2144] = 6'b111110;
		color_arr[2145] = 6'b111110;
		color_arr[2146] = 6'b111110;
		color_arr[2147] = 6'b111110;
		color_arr[2148] = 6'b111010;
		color_arr[2149] = 6'b111010;
		color_arr[2150] = 6'b111001;
		color_arr[2151] = 6'b111001;
		color_arr[2152] = 6'b111001;
		color_arr[2153] = 6'b111001;
		color_arr[2154] = 6'b111001;
		color_arr[2155] = 6'b111010;
		color_arr[2156] = 6'b111110;
		color_arr[2157] = 6'b111001;
		color_arr[2158] = 6'b111001;
		color_arr[2159] = 6'b000000;
		color_arr[2160] = 6'b000000;
		color_arr[2161] = 6'b000000;
		color_arr[2162] = 6'b000000;
		color_arr[2163] = 6'b000000;
		color_arr[2164] = 6'b000000;
		color_arr[2165] = 6'b000000;
		color_arr[2166] = 6'b000000;
		color_arr[2167] = 6'b000000;
		color_arr[2168] = 6'b000000;
		color_arr[2169] = 6'b000000;
		color_arr[2170] = 6'b000000;
		color_arr[2171] = 6'b000000;
		color_arr[2172] = 6'b000000;
		color_arr[2173] = 6'b000000;
		color_arr[2174] = 6'b000000;
		color_arr[2175] = 6'b000000;
		color_arr[2176] = 6'b000000;
		color_arr[2177] = 6'b000000;
		color_arr[2178] = 6'b000000;
		color_arr[2179] = 6'b000000;
		color_arr[2180] = 6'b000000;
		color_arr[2181] = 6'b000000;
		color_arr[2182] = 6'b000000;
		color_arr[2183] = 6'b000000;
		color_arr[2184] = 6'b000000;
		color_arr[2185] = 6'b000000;
		color_arr[2186] = 6'b000000;
		color_arr[2187] = 6'b000000;
		color_arr[2188] = 6'b000000;
		color_arr[2189] = 6'b000000;
		color_arr[2190] = 6'b000000;
		color_arr[2191] = 6'b000000;
		color_arr[2192] = 6'b000000;
		color_arr[2193] = 6'b000000;
		color_arr[2194] = 6'b000000;
		color_arr[2195] = 6'b000000;
		color_arr[2196] = 6'b111110;
		color_arr[2197] = 6'b111110;
		color_arr[2198] = 6'b111110;
		color_arr[2199] = 6'b111110;
		color_arr[2200] = 6'b111110;
		color_arr[2201] = 6'b111110;
		color_arr[2202] = 6'b111110;
		color_arr[2203] = 6'b111110;
		color_arr[2204] = 6'b111110;
		color_arr[2205] = 6'b111110;
		color_arr[2206] = 6'b111110;
		color_arr[2207] = 6'b111110;
		color_arr[2208] = 6'b111110;
		color_arr[2209] = 6'b111110;
		color_arr[2210] = 6'b111110;
		color_arr[2211] = 6'b111110;
		color_arr[2212] = 6'b111110;
		color_arr[2213] = 6'b111001;
		color_arr[2214] = 6'b111001;
		color_arr[2215] = 6'b111001;
		color_arr[2216] = 6'b111001;
		color_arr[2217] = 6'b111001;
		color_arr[2218] = 6'b111010;
		color_arr[2219] = 6'b111110;
		color_arr[2220] = 6'b111110;
		color_arr[2221] = 6'b111110;
		color_arr[2222] = 6'b111001;
		color_arr[2223] = 6'b111001;
		color_arr[2224] = 6'b000000;
		color_arr[2225] = 6'b000000;
		color_arr[2226] = 6'b000000;
		color_arr[2227] = 6'b000000;
		color_arr[2228] = 6'b000000;
		color_arr[2229] = 6'b000000;
		color_arr[2230] = 6'b000000;
		color_arr[2231] = 6'b000000;
		color_arr[2232] = 6'b000000;
		color_arr[2233] = 6'b000000;
		color_arr[2234] = 6'b000000;
		color_arr[2235] = 6'b000000;
		color_arr[2236] = 6'b000000;
		color_arr[2237] = 6'b000000;
		color_arr[2238] = 6'b000000;
		color_arr[2239] = 6'b000000;
		color_arr[2240] = 6'b000000;
		color_arr[2241] = 6'b000000;
		color_arr[2242] = 6'b000000;
		color_arr[2243] = 6'b000000;
		color_arr[2244] = 6'b000000;
		color_arr[2245] = 6'b000000;
		color_arr[2246] = 6'b000000;
		color_arr[2247] = 6'b000000;
		color_arr[2248] = 6'b000000;
		color_arr[2249] = 6'b000000;
		color_arr[2250] = 6'b000000;
		color_arr[2251] = 6'b000000;
		color_arr[2252] = 6'b000000;
		color_arr[2253] = 6'b000000;
		color_arr[2254] = 6'b000000;
		color_arr[2255] = 6'b000000;
		color_arr[2256] = 6'b000000;
		color_arr[2257] = 6'b000000;
		color_arr[2258] = 6'b000000;
		color_arr[2259] = 6'b111110;
		color_arr[2260] = 6'b111110;
		color_arr[2261] = 6'b111110;
		color_arr[2262] = 6'b111110;
		color_arr[2263] = 6'b111110;
		color_arr[2264] = 6'b111110;
		color_arr[2265] = 6'b111110;
		color_arr[2266] = 6'b111110;
		color_arr[2267] = 6'b111110;
		color_arr[2268] = 6'b111110;
		color_arr[2269] = 6'b111110;
		color_arr[2270] = 6'b111110;
		color_arr[2271] = 6'b111110;
		color_arr[2272] = 6'b111110;
		color_arr[2273] = 6'b111110;
		color_arr[2274] = 6'b111110;
		color_arr[2275] = 6'b111110;
		color_arr[2276] = 6'b111110;
		color_arr[2277] = 6'b111010;
		color_arr[2278] = 6'b111001;
		color_arr[2279] = 6'b111010;
		color_arr[2280] = 6'b111010;
		color_arr[2281] = 6'b111110;
		color_arr[2282] = 6'b111110;
		color_arr[2283] = 6'b111110;
		color_arr[2284] = 6'b111110;
		color_arr[2285] = 6'b111110;
		color_arr[2286] = 6'b111110;
		color_arr[2287] = 6'b111001;
		color_arr[2288] = 6'b000000;
		color_arr[2289] = 6'b000000;
		color_arr[2290] = 6'b000000;
		color_arr[2291] = 6'b000000;
		color_arr[2292] = 6'b000000;
		color_arr[2293] = 6'b000000;
		color_arr[2294] = 6'b000000;
		color_arr[2295] = 6'b000000;
		color_arr[2296] = 6'b000000;
		color_arr[2297] = 6'b000000;
		color_arr[2298] = 6'b000000;
		color_arr[2299] = 6'b000000;
		color_arr[2300] = 6'b000000;
		color_arr[2301] = 6'b000000;
		color_arr[2302] = 6'b000000;
		color_arr[2303] = 6'b000000;
		color_arr[2304] = 6'b000000;
		color_arr[2305] = 6'b000000;
		color_arr[2306] = 6'b000000;
		color_arr[2307] = 6'b000000;
		color_arr[2308] = 6'b000000;
		color_arr[2309] = 6'b000000;
		color_arr[2310] = 6'b000000;
		color_arr[2311] = 6'b000000;
		color_arr[2312] = 6'b000000;
		color_arr[2313] = 6'b000000;
		color_arr[2314] = 6'b000000;
		color_arr[2315] = 6'b000000;
		color_arr[2316] = 6'b000000;
		color_arr[2317] = 6'b000000;
		color_arr[2318] = 6'b000000;
		color_arr[2319] = 6'b000000;
		color_arr[2320] = 6'b000000;
		color_arr[2321] = 6'b000000;
		color_arr[2322] = 6'b000000;
		color_arr[2323] = 6'b111110;
		color_arr[2324] = 6'b111110;
		color_arr[2325] = 6'b111110;
		color_arr[2326] = 6'b111110;
		color_arr[2327] = 6'b111110;
		color_arr[2328] = 6'b111110;
		color_arr[2329] = 6'b111110;
		color_arr[2330] = 6'b111110;
		color_arr[2331] = 6'b111110;
		color_arr[2332] = 6'b111110;
		color_arr[2333] = 6'b111110;
		color_arr[2334] = 6'b111110;
		color_arr[2335] = 6'b111110;
		color_arr[2336] = 6'b111110;
		color_arr[2337] = 6'b111110;
		color_arr[2338] = 6'b111110;
		color_arr[2339] = 6'b111110;
		color_arr[2340] = 6'b111110;
		color_arr[2341] = 6'b111110;
		color_arr[2342] = 6'b111110;
		color_arr[2343] = 6'b111110;
		color_arr[2344] = 6'b111110;
		color_arr[2345] = 6'b111110;
		color_arr[2346] = 6'b111110;
		color_arr[2347] = 6'b111110;
		color_arr[2348] = 6'b111110;
		color_arr[2349] = 6'b111110;
		color_arr[2350] = 6'b111110;
		color_arr[2351] = 6'b111001;
		color_arr[2352] = 6'b000000;
		color_arr[2353] = 6'b000000;
		color_arr[2354] = 6'b000000;
		color_arr[2355] = 6'b000000;
		color_arr[2356] = 6'b000000;
		color_arr[2357] = 6'b000000;
		color_arr[2358] = 6'b000000;
		color_arr[2359] = 6'b000000;
		color_arr[2360] = 6'b000000;
		color_arr[2361] = 6'b000000;
		color_arr[2362] = 6'b000000;
		color_arr[2363] = 6'b000000;
		color_arr[2364] = 6'b000000;
		color_arr[2365] = 6'b000000;
		color_arr[2366] = 6'b000000;
		color_arr[2367] = 6'b000000;
		color_arr[2368] = 6'b000000;
		color_arr[2369] = 6'b000000;
		color_arr[2370] = 6'b000000;
		color_arr[2371] = 6'b000000;
		color_arr[2372] = 6'b000000;
		color_arr[2373] = 6'b000000;
		color_arr[2374] = 6'b000000;
		color_arr[2375] = 6'b000000;
		color_arr[2376] = 6'b000000;
		color_arr[2377] = 6'b000000;
		color_arr[2378] = 6'b000000;
		color_arr[2379] = 6'b000000;
		color_arr[2380] = 6'b000000;
		color_arr[2381] = 6'b000000;
		color_arr[2382] = 6'b000000;
		color_arr[2383] = 6'b000000;
		color_arr[2384] = 6'b000000;
		color_arr[2385] = 6'b000000;
		color_arr[2386] = 6'b111110;
		color_arr[2387] = 6'b111110;
		color_arr[2388] = 6'b111110;
		color_arr[2389] = 6'b111110;
		color_arr[2390] = 6'b111110;
		color_arr[2391] = 6'b111110;
		color_arr[2392] = 6'b111110;
		color_arr[2393] = 6'b111110;
		color_arr[2394] = 6'b111110;
		color_arr[2395] = 6'b111110;
		color_arr[2396] = 6'b111110;
		color_arr[2397] = 6'b111110;
		color_arr[2398] = 6'b111110;
		color_arr[2399] = 6'b111110;
		color_arr[2400] = 6'b111110;
		color_arr[2401] = 6'b111110;
		color_arr[2402] = 6'b111110;
		color_arr[2403] = 6'b111110;
		color_arr[2404] = 6'b111110;
		color_arr[2405] = 6'b111110;
		color_arr[2406] = 6'b111110;
		color_arr[2407] = 6'b111110;
		color_arr[2408] = 6'b111110;
		color_arr[2409] = 6'b111110;
		color_arr[2410] = 6'b111110;
		color_arr[2411] = 6'b111110;
		color_arr[2412] = 6'b111110;
		color_arr[2413] = 6'b111110;
		color_arr[2414] = 6'b111110;
		color_arr[2415] = 6'b111001;
		color_arr[2416] = 6'b000000;
		color_arr[2417] = 6'b000000;
		color_arr[2418] = 6'b000000;
		color_arr[2419] = 6'b000000;
		color_arr[2420] = 6'b000000;
		color_arr[2421] = 6'b000000;
		color_arr[2422] = 6'b000000;
		color_arr[2423] = 6'b000000;
		color_arr[2424] = 6'b000000;
		color_arr[2425] = 6'b000000;
		color_arr[2426] = 6'b000000;
		color_arr[2427] = 6'b000000;
		color_arr[2428] = 6'b000000;
		color_arr[2429] = 6'b000000;
		color_arr[2430] = 6'b000000;
		color_arr[2431] = 6'b000000;
		color_arr[2432] = 6'b000000;
		color_arr[2433] = 6'b000000;
		color_arr[2434] = 6'b000000;
		color_arr[2435] = 6'b000000;
		color_arr[2436] = 6'b000000;
		color_arr[2437] = 6'b000000;
		color_arr[2438] = 6'b000000;
		color_arr[2439] = 6'b000000;
		color_arr[2440] = 6'b000000;
		color_arr[2441] = 6'b000000;
		color_arr[2442] = 6'b000000;
		color_arr[2443] = 6'b000000;
		color_arr[2444] = 6'b000000;
		color_arr[2445] = 6'b000000;
		color_arr[2446] = 6'b000000;
		color_arr[2447] = 6'b000000;
		color_arr[2448] = 6'b000000;
		color_arr[2449] = 6'b000000;
		color_arr[2450] = 6'b111110;
		color_arr[2451] = 6'b111110;
		color_arr[2452] = 6'b111110;
		color_arr[2453] = 6'b111110;
		color_arr[2454] = 6'b111110;
		color_arr[2455] = 6'b111110;
		color_arr[2456] = 6'b111110;
		color_arr[2457] = 6'b111110;
		color_arr[2458] = 6'b111110;
		color_arr[2459] = 6'b111110;
		color_arr[2460] = 6'b111110;
		color_arr[2461] = 6'b111110;
		color_arr[2462] = 6'b111110;
		color_arr[2463] = 6'b111110;
		color_arr[2464] = 6'b111110;
		color_arr[2465] = 6'b111110;
		color_arr[2466] = 6'b111110;
		color_arr[2467] = 6'b111110;
		color_arr[2468] = 6'b111110;
		color_arr[2469] = 6'b111110;
		color_arr[2470] = 6'b111110;
		color_arr[2471] = 6'b111110;
		color_arr[2472] = 6'b111110;
		color_arr[2473] = 6'b111110;
		color_arr[2474] = 6'b111110;
		color_arr[2475] = 6'b111110;
		color_arr[2476] = 6'b111110;
		color_arr[2477] = 6'b111110;
		color_arr[2478] = 6'b111110;
		color_arr[2479] = 6'b111001;
		color_arr[2480] = 6'b111001;
		color_arr[2481] = 6'b000000;
		color_arr[2482] = 6'b000000;
		color_arr[2483] = 6'b000000;
		color_arr[2484] = 6'b000000;
		color_arr[2485] = 6'b000000;
		color_arr[2486] = 6'b000000;
		color_arr[2487] = 6'b000000;
		color_arr[2488] = 6'b000000;
		color_arr[2489] = 6'b000000;
		color_arr[2490] = 6'b000000;
		color_arr[2491] = 6'b000000;
		color_arr[2492] = 6'b000000;
		color_arr[2493] = 6'b000000;
		color_arr[2494] = 6'b000000;
		color_arr[2495] = 6'b000000;
		color_arr[2496] = 6'b000000;
		color_arr[2497] = 6'b000000;
		color_arr[2498] = 6'b000000;
		color_arr[2499] = 6'b000000;
		color_arr[2500] = 6'b000000;
		color_arr[2501] = 6'b000000;
		color_arr[2502] = 6'b000000;
		color_arr[2503] = 6'b000000;
		color_arr[2504] = 6'b000000;
		color_arr[2505] = 6'b000000;
		color_arr[2506] = 6'b000000;
		color_arr[2507] = 6'b000000;
		color_arr[2508] = 6'b000000;
		color_arr[2509] = 6'b000000;
		color_arr[2510] = 6'b000000;
		color_arr[2511] = 6'b000000;
		color_arr[2512] = 6'b000000;
		color_arr[2513] = 6'b000000;
		color_arr[2514] = 6'b111110;
		color_arr[2515] = 6'b111110;
		color_arr[2516] = 6'b111110;
		color_arr[2517] = 6'b111110;
		color_arr[2518] = 6'b111110;
		color_arr[2519] = 6'b111110;
		color_arr[2520] = 6'b111110;
		color_arr[2521] = 6'b111110;
		color_arr[2522] = 6'b111110;
		color_arr[2523] = 6'b111110;
		color_arr[2524] = 6'b111110;
		color_arr[2525] = 6'b111110;
		color_arr[2526] = 6'b111110;
		color_arr[2527] = 6'b111110;
		color_arr[2528] = 6'b111110;
		color_arr[2529] = 6'b111110;
		color_arr[2530] = 6'b111110;
		color_arr[2531] = 6'b111110;
		color_arr[2532] = 6'b111110;
		color_arr[2533] = 6'b111110;
		color_arr[2534] = 6'b111110;
		color_arr[2535] = 6'b111110;
		color_arr[2536] = 6'b111110;
		color_arr[2537] = 6'b111110;
		color_arr[2538] = 6'b111110;
		color_arr[2539] = 6'b111110;
		color_arr[2540] = 6'b111110;
		color_arr[2541] = 6'b111110;
		color_arr[2542] = 6'b111010;
		color_arr[2543] = 6'b111001;
		color_arr[2544] = 6'b111001;
		color_arr[2545] = 6'b000000;
		color_arr[2546] = 6'b000000;
		color_arr[2547] = 6'b000000;
		color_arr[2548] = 6'b000000;
		color_arr[2549] = 6'b000000;
		color_arr[2550] = 6'b000000;
		color_arr[2551] = 6'b000000;
		color_arr[2552] = 6'b000000;
		color_arr[2553] = 6'b000000;
		color_arr[2554] = 6'b000000;
		color_arr[2555] = 6'b000000;
		color_arr[2556] = 6'b000000;
		color_arr[2557] = 6'b000000;
		color_arr[2558] = 6'b000000;
		color_arr[2559] = 6'b000000;
		color_arr[2560] = 6'b000000;
		color_arr[2561] = 6'b000000;
		color_arr[2562] = 6'b000000;
		color_arr[2563] = 6'b000000;
		color_arr[2564] = 6'b000000;
		color_arr[2565] = 6'b000000;
		color_arr[2566] = 6'b000000;
		color_arr[2567] = 6'b000000;
		color_arr[2568] = 6'b000000;
		color_arr[2569] = 6'b000000;
		color_arr[2570] = 6'b000000;
		color_arr[2571] = 6'b000000;
		color_arr[2572] = 6'b000000;
		color_arr[2573] = 6'b000000;
		color_arr[2574] = 6'b000000;
		color_arr[2575] = 6'b000000;
		color_arr[2576] = 6'b000000;
		color_arr[2577] = 6'b111110;
		color_arr[2578] = 6'b111110;
		color_arr[2579] = 6'b111110;
		color_arr[2580] = 6'b111110;
		color_arr[2581] = 6'b111110;
		color_arr[2582] = 6'b111110;
		color_arr[2583] = 6'b111110;
		color_arr[2584] = 6'b111110;
		color_arr[2585] = 6'b111110;
		color_arr[2586] = 6'b111110;
		color_arr[2587] = 6'b111110;
		color_arr[2588] = 6'b111110;
		color_arr[2589] = 6'b111110;
		color_arr[2590] = 6'b111110;
		color_arr[2591] = 6'b111110;
		color_arr[2592] = 6'b111110;
		color_arr[2593] = 6'b111110;
		color_arr[2594] = 6'b111110;
		color_arr[2595] = 6'b111110;
		color_arr[2596] = 6'b111110;
		color_arr[2597] = 6'b111110;
		color_arr[2598] = 6'b111110;
		color_arr[2599] = 6'b111110;
		color_arr[2600] = 6'b111110;
		color_arr[2601] = 6'b111110;
		color_arr[2602] = 6'b111110;
		color_arr[2603] = 6'b111110;
		color_arr[2604] = 6'b111110;
		color_arr[2605] = 6'b111010;
		color_arr[2606] = 6'b111001;
		color_arr[2607] = 6'b111001;
		color_arr[2608] = 6'b111001;
		color_arr[2609] = 6'b000000;
		color_arr[2610] = 6'b000000;
		color_arr[2611] = 6'b000000;
		color_arr[2612] = 6'b000000;
		color_arr[2613] = 6'b000000;
		color_arr[2614] = 6'b000000;
		color_arr[2615] = 6'b000000;
		color_arr[2616] = 6'b000000;
		color_arr[2617] = 6'b000000;
		color_arr[2618] = 6'b000000;
		color_arr[2619] = 6'b000000;
		color_arr[2620] = 6'b000000;
		color_arr[2621] = 6'b000000;
		color_arr[2622] = 6'b000000;
		color_arr[2623] = 6'b000000;
		color_arr[2624] = 6'b000000;
		color_arr[2625] = 6'b000000;
		color_arr[2626] = 6'b000000;
		color_arr[2627] = 6'b000000;
		color_arr[2628] = 6'b000000;
		color_arr[2629] = 6'b000000;
		color_arr[2630] = 6'b000000;
		color_arr[2631] = 6'b000000;
		color_arr[2632] = 6'b000000;
		color_arr[2633] = 6'b000000;
		color_arr[2634] = 6'b000000;
		color_arr[2635] = 6'b000000;
		color_arr[2636] = 6'b000000;
		color_arr[2637] = 6'b000000;
		color_arr[2638] = 6'b000000;
		color_arr[2639] = 6'b000000;
		color_arr[2640] = 6'b000000;
		color_arr[2641] = 6'b111110;
		color_arr[2642] = 6'b111110;
		color_arr[2643] = 6'b111110;
		color_arr[2644] = 6'b111110;
		color_arr[2645] = 6'b111110;
		color_arr[2646] = 6'b111110;
		color_arr[2647] = 6'b111110;
		color_arr[2648] = 6'b111110;
		color_arr[2649] = 6'b111110;
		color_arr[2650] = 6'b111110;
		color_arr[2651] = 6'b111110;
		color_arr[2652] = 6'b111110;
		color_arr[2653] = 6'b111110;
		color_arr[2654] = 6'b111110;
		color_arr[2655] = 6'b111110;
		color_arr[2656] = 6'b111110;
		color_arr[2657] = 6'b111110;
		color_arr[2658] = 6'b111110;
		color_arr[2659] = 6'b111110;
		color_arr[2660] = 6'b111110;
		color_arr[2661] = 6'b111110;
		color_arr[2662] = 6'b111110;
		color_arr[2663] = 6'b111110;
		color_arr[2664] = 6'b111110;
		color_arr[2665] = 6'b111110;
		color_arr[2666] = 6'b111110;
		color_arr[2667] = 6'b111110;
		color_arr[2668] = 6'b111010;
		color_arr[2669] = 6'b111001;
		color_arr[2670] = 6'b111001;
		color_arr[2671] = 6'b111001;
		color_arr[2672] = 6'b111001;
		color_arr[2673] = 6'b000000;
		color_arr[2674] = 6'b000000;
		color_arr[2675] = 6'b000000;
		color_arr[2676] = 6'b000000;
		color_arr[2677] = 6'b000000;
		color_arr[2678] = 6'b000000;
		color_arr[2679] = 6'b000000;
		color_arr[2680] = 6'b000000;
		color_arr[2681] = 6'b000000;
		color_arr[2682] = 6'b000000;
		color_arr[2683] = 6'b000000;
		color_arr[2684] = 6'b000000;
		color_arr[2685] = 6'b000000;
		color_arr[2686] = 6'b000000;
		color_arr[2687] = 6'b000000;
		color_arr[2688] = 6'b000000;
		color_arr[2689] = 6'b000000;
		color_arr[2690] = 6'b000000;
		color_arr[2691] = 6'b000000;
		color_arr[2692] = 6'b000000;
		color_arr[2693] = 6'b000000;
		color_arr[2694] = 6'b000000;
		color_arr[2695] = 6'b000000;
		color_arr[2696] = 6'b000000;
		color_arr[2697] = 6'b000000;
		color_arr[2698] = 6'b000000;
		color_arr[2699] = 6'b000000;
		color_arr[2700] = 6'b000000;
		color_arr[2701] = 6'b000000;
		color_arr[2702] = 6'b000000;
		color_arr[2703] = 6'b000000;
		color_arr[2704] = 6'b111110;
		color_arr[2705] = 6'b111110;
		color_arr[2706] = 6'b111110;
		color_arr[2707] = 6'b111110;
		color_arr[2708] = 6'b111110;
		color_arr[2709] = 6'b111110;
		color_arr[2710] = 6'b111110;
		color_arr[2711] = 6'b111110;
		color_arr[2712] = 6'b111110;
		color_arr[2713] = 6'b111110;
		color_arr[2714] = 6'b111110;
		color_arr[2715] = 6'b111110;
		color_arr[2716] = 6'b111110;
		color_arr[2717] = 6'b111110;
		color_arr[2718] = 6'b111110;
		color_arr[2719] = 6'b111110;
		color_arr[2720] = 6'b111110;
		color_arr[2721] = 6'b111110;
		color_arr[2722] = 6'b111110;
		color_arr[2723] = 6'b111110;
		color_arr[2724] = 6'b111110;
		color_arr[2725] = 6'b111110;
		color_arr[2726] = 6'b111110;
		color_arr[2727] = 6'b111110;
		color_arr[2728] = 6'b111110;
		color_arr[2729] = 6'b111110;
		color_arr[2730] = 6'b111110;
		color_arr[2731] = 6'b111110;
		color_arr[2732] = 6'b111110;
		color_arr[2733] = 6'b111110;
		color_arr[2734] = 6'b111010;
		color_arr[2735] = 6'b111001;
		color_arr[2736] = 6'b111001;
		color_arr[2737] = 6'b000000;
		color_arr[2738] = 6'b000000;
		color_arr[2739] = 6'b000000;
		color_arr[2740] = 6'b000000;
		color_arr[2741] = 6'b000000;
		color_arr[2742] = 6'b000000;
		color_arr[2743] = 6'b000000;
		color_arr[2744] = 6'b000000;
		color_arr[2745] = 6'b000000;
		color_arr[2746] = 6'b000000;
		color_arr[2747] = 6'b000000;
		color_arr[2748] = 6'b000000;
		color_arr[2749] = 6'b000000;
		color_arr[2750] = 6'b000000;
		color_arr[2751] = 6'b000000;
		color_arr[2752] = 6'b000000;
		color_arr[2753] = 6'b000000;
		color_arr[2754] = 6'b000000;
		color_arr[2755] = 6'b000000;
		color_arr[2756] = 6'b000000;
		color_arr[2757] = 6'b000000;
		color_arr[2758] = 6'b000000;
		color_arr[2759] = 6'b000000;
		color_arr[2760] = 6'b000000;
		color_arr[2761] = 6'b000000;
		color_arr[2762] = 6'b000000;
		color_arr[2763] = 6'b000000;
		color_arr[2764] = 6'b000000;
		color_arr[2765] = 6'b000000;
		color_arr[2766] = 6'b000000;
		color_arr[2767] = 6'b000000;
		color_arr[2768] = 6'b111010;
		color_arr[2769] = 6'b111110;
		color_arr[2770] = 6'b111110;
		color_arr[2771] = 6'b111110;
		color_arr[2772] = 6'b111110;
		color_arr[2773] = 6'b111110;
		color_arr[2774] = 6'b111110;
		color_arr[2775] = 6'b111110;
		color_arr[2776] = 6'b111110;
		color_arr[2777] = 6'b111110;
		color_arr[2778] = 6'b111110;
		color_arr[2779] = 6'b111110;
		color_arr[2780] = 6'b111110;
		color_arr[2781] = 6'b111110;
		color_arr[2782] = 6'b111110;
		color_arr[2783] = 6'b111110;
		color_arr[2784] = 6'b111110;
		color_arr[2785] = 6'b111110;
		color_arr[2786] = 6'b111110;
		color_arr[2787] = 6'b111110;
		color_arr[2788] = 6'b111110;
		color_arr[2789] = 6'b111110;
		color_arr[2790] = 6'b111110;
		color_arr[2791] = 6'b111110;
		color_arr[2792] = 6'b111110;
		color_arr[2793] = 6'b111110;
		color_arr[2794] = 6'b111110;
		color_arr[2795] = 6'b111110;
		color_arr[2796] = 6'b111110;
		color_arr[2797] = 6'b111110;
		color_arr[2798] = 6'b111110;
		color_arr[2799] = 6'b111010;
		color_arr[2800] = 6'b111001;
		color_arr[2801] = 6'b000000;
		color_arr[2802] = 6'b000000;
		color_arr[2803] = 6'b000000;
		color_arr[2804] = 6'b000000;
		color_arr[2805] = 6'b000000;
		color_arr[2806] = 6'b000000;
		color_arr[2807] = 6'b000000;
		color_arr[2808] = 6'b000000;
		color_arr[2809] = 6'b000000;
		color_arr[2810] = 6'b000000;
		color_arr[2811] = 6'b000000;
		color_arr[2812] = 6'b000000;
		color_arr[2813] = 6'b000000;
		color_arr[2814] = 6'b000000;
		color_arr[2815] = 6'b000000;
		color_arr[2816] = 6'b000000;
		color_arr[2817] = 6'b000000;
		color_arr[2818] = 6'b000000;
		color_arr[2819] = 6'b000000;
		color_arr[2820] = 6'b000000;
		color_arr[2821] = 6'b000000;
		color_arr[2822] = 6'b000000;
		color_arr[2823] = 6'b000000;
		color_arr[2824] = 6'b000000;
		color_arr[2825] = 6'b000000;
		color_arr[2826] = 6'b000000;
		color_arr[2827] = 6'b000000;
		color_arr[2828] = 6'b000000;
		color_arr[2829] = 6'b000000;
		color_arr[2830] = 6'b000000;
		color_arr[2831] = 6'b000000;
		color_arr[2832] = 6'b111001;
		color_arr[2833] = 6'b111110;
		color_arr[2834] = 6'b111110;
		color_arr[2835] = 6'b111110;
		color_arr[2836] = 6'b111110;
		color_arr[2837] = 6'b111110;
		color_arr[2838] = 6'b111110;
		color_arr[2839] = 6'b111110;
		color_arr[2840] = 6'b111110;
		color_arr[2841] = 6'b111110;
		color_arr[2842] = 6'b111110;
		color_arr[2843] = 6'b111110;
		color_arr[2844] = 6'b111110;
		color_arr[2845] = 6'b111110;
		color_arr[2846] = 6'b111110;
		color_arr[2847] = 6'b111110;
		color_arr[2848] = 6'b111110;
		color_arr[2849] = 6'b111110;
		color_arr[2850] = 6'b111110;
		color_arr[2851] = 6'b111110;
		color_arr[2852] = 6'b111110;
		color_arr[2853] = 6'b111110;
		color_arr[2854] = 6'b111110;
		color_arr[2855] = 6'b111110;
		color_arr[2856] = 6'b111110;
		color_arr[2857] = 6'b111110;
		color_arr[2858] = 6'b111110;
		color_arr[2859] = 6'b111110;
		color_arr[2860] = 6'b111110;
		color_arr[2861] = 6'b111110;
		color_arr[2862] = 6'b111110;
		color_arr[2863] = 6'b111010;
		color_arr[2864] = 6'b111001;
		color_arr[2865] = 6'b000000;
		color_arr[2866] = 6'b000000;
		color_arr[2867] = 6'b000000;
		color_arr[2868] = 6'b000000;
		color_arr[2869] = 6'b000000;
		color_arr[2870] = 6'b000000;
		color_arr[2871] = 6'b000000;
		color_arr[2872] = 6'b000000;
		color_arr[2873] = 6'b000000;
		color_arr[2874] = 6'b000000;
		color_arr[2875] = 6'b000000;
		color_arr[2876] = 6'b000000;
		color_arr[2877] = 6'b000000;
		color_arr[2878] = 6'b000000;
		color_arr[2879] = 6'b000000;
		color_arr[2880] = 6'b000000;
		color_arr[2881] = 6'b000000;
		color_arr[2882] = 6'b000000;
		color_arr[2883] = 6'b000000;
		color_arr[2884] = 6'b000000;
		color_arr[2885] = 6'b000000;
		color_arr[2886] = 6'b000000;
		color_arr[2887] = 6'b000000;
		color_arr[2888] = 6'b000000;
		color_arr[2889] = 6'b000000;
		color_arr[2890] = 6'b000000;
		color_arr[2891] = 6'b000000;
		color_arr[2892] = 6'b000000;
		color_arr[2893] = 6'b000000;
		color_arr[2894] = 6'b000000;
		color_arr[2895] = 6'b111001;
		color_arr[2896] = 6'b111010;
		color_arr[2897] = 6'b111110;
		color_arr[2898] = 6'b111110;
		color_arr[2899] = 6'b111110;
		color_arr[2900] = 6'b111110;
		color_arr[2901] = 6'b111110;
		color_arr[2902] = 6'b111110;
		color_arr[2903] = 6'b111110;
		color_arr[2904] = 6'b111110;
		color_arr[2905] = 6'b111110;
		color_arr[2906] = 6'b111110;
		color_arr[2907] = 6'b111110;
		color_arr[2908] = 6'b111110;
		color_arr[2909] = 6'b111110;
		color_arr[2910] = 6'b111110;
		color_arr[2911] = 6'b111110;
		color_arr[2912] = 6'b111110;
		color_arr[2913] = 6'b111110;
		color_arr[2914] = 6'b111110;
		color_arr[2915] = 6'b111110;
		color_arr[2916] = 6'b111110;
		color_arr[2917] = 6'b111110;
		color_arr[2918] = 6'b111110;
		color_arr[2919] = 6'b111110;
		color_arr[2920] = 6'b111110;
		color_arr[2921] = 6'b111110;
		color_arr[2922] = 6'b111110;
		color_arr[2923] = 6'b111110;
		color_arr[2924] = 6'b111110;
		color_arr[2925] = 6'b111110;
		color_arr[2926] = 6'b111110;
		color_arr[2927] = 6'b111110;
		color_arr[2928] = 6'b111001;
		color_arr[2929] = 6'b000000;
		color_arr[2930] = 6'b000000;
		color_arr[2931] = 6'b000000;
		color_arr[2932] = 6'b000000;
		color_arr[2933] = 6'b000000;
		color_arr[2934] = 6'b000000;
		color_arr[2935] = 6'b000000;
		color_arr[2936] = 6'b000000;
		color_arr[2937] = 6'b000000;
		color_arr[2938] = 6'b000000;
		color_arr[2939] = 6'b000000;
		color_arr[2940] = 6'b000000;
		color_arr[2941] = 6'b000000;
		color_arr[2942] = 6'b000000;
		color_arr[2943] = 6'b000000;
		color_arr[2944] = 6'b000000;
		color_arr[2945] = 6'b000000;
		color_arr[2946] = 6'b000000;
		color_arr[2947] = 6'b000000;
		color_arr[2948] = 6'b000000;
		color_arr[2949] = 6'b000000;
		color_arr[2950] = 6'b000000;
		color_arr[2951] = 6'b000000;
		color_arr[2952] = 6'b000000;
		color_arr[2953] = 6'b000000;
		color_arr[2954] = 6'b000000;
		color_arr[2955] = 6'b000000;
		color_arr[2956] = 6'b000000;
		color_arr[2957] = 6'b000000;
		color_arr[2958] = 6'b000000;
		color_arr[2959] = 6'b111001;
		color_arr[2960] = 6'b111010;
		color_arr[2961] = 6'b111010;
		color_arr[2962] = 6'b111010;
		color_arr[2963] = 6'b111010;
		color_arr[2964] = 6'b111010;
		color_arr[2965] = 6'b111110;
		color_arr[2966] = 6'b111110;
		color_arr[2967] = 6'b111001;
		color_arr[2968] = 6'b111001;
		color_arr[2969] = 6'b111110;
		color_arr[2970] = 6'b111110;
		color_arr[2971] = 6'b111110;
		color_arr[2972] = 6'b111110;
		color_arr[2973] = 6'b111110;
		color_arr[2974] = 6'b111110;
		color_arr[2975] = 6'b111110;
		color_arr[2976] = 6'b111110;
		color_arr[2977] = 6'b111110;
		color_arr[2978] = 6'b111110;
		color_arr[2979] = 6'b111110;
		color_arr[2980] = 6'b111110;
		color_arr[2981] = 6'b111110;
		color_arr[2982] = 6'b111110;
		color_arr[2983] = 6'b111110;
		color_arr[2984] = 6'b111110;
		color_arr[2985] = 6'b111110;
		color_arr[2986] = 6'b111110;
		color_arr[2987] = 6'b111110;
		color_arr[2988] = 6'b111110;
		color_arr[2989] = 6'b111110;
		color_arr[2990] = 6'b111110;
		color_arr[2991] = 6'b111110;
		color_arr[2992] = 6'b111001;
		color_arr[2993] = 6'b000000;
		color_arr[2994] = 6'b000000;
		color_arr[2995] = 6'b000000;
		color_arr[2996] = 6'b000000;
		color_arr[2997] = 6'b000000;
		color_arr[2998] = 6'b000000;
		color_arr[2999] = 6'b000000;
		color_arr[3000] = 6'b000000;
		color_arr[3001] = 6'b000000;
		color_arr[3002] = 6'b000000;
		color_arr[3003] = 6'b000000;
		color_arr[3004] = 6'b000000;
		color_arr[3005] = 6'b000000;
		color_arr[3006] = 6'b000000;
		color_arr[3007] = 6'b000000;
		color_arr[3008] = 6'b000000;
		color_arr[3009] = 6'b000000;
		color_arr[3010] = 6'b000000;
		color_arr[3011] = 6'b000000;
		color_arr[3012] = 6'b000000;
		color_arr[3013] = 6'b000000;
		color_arr[3014] = 6'b000000;
		color_arr[3015] = 6'b000000;
		color_arr[3016] = 6'b000000;
		color_arr[3017] = 6'b000000;
		color_arr[3018] = 6'b000000;
		color_arr[3019] = 6'b000000;
		color_arr[3020] = 6'b000000;
		color_arr[3021] = 6'b000000;
		color_arr[3022] = 6'b000000;
		color_arr[3023] = 6'b111001;
		color_arr[3024] = 6'b111001;
		color_arr[3025] = 6'b111010;
		color_arr[3026] = 6'b111010;
		color_arr[3027] = 6'b111010;
		color_arr[3028] = 6'b111010;
		color_arr[3029] = 6'b111010;
		color_arr[3030] = 6'b111010;
		color_arr[3031] = 6'b111010;
		color_arr[3032] = 6'b111010;
		color_arr[3033] = 6'b111001;
		color_arr[3034] = 6'b111001;
		color_arr[3035] = 6'b111110;
		color_arr[3036] = 6'b111110;
		color_arr[3037] = 6'b111110;
		color_arr[3038] = 6'b111010;
		color_arr[3039] = 6'b111001;
		color_arr[3040] = 6'b111001;
		color_arr[3041] = 6'b111001;
		color_arr[3042] = 6'b111110;
		color_arr[3043] = 6'b111110;
		color_arr[3044] = 6'b111110;
		color_arr[3045] = 6'b111110;
		color_arr[3046] = 6'b111110;
		color_arr[3047] = 6'b111110;
		color_arr[3048] = 6'b111110;
		color_arr[3049] = 6'b111110;
		color_arr[3050] = 6'b111110;
		color_arr[3051] = 6'b111110;
		color_arr[3052] = 6'b111110;
		color_arr[3053] = 6'b111010;
		color_arr[3054] = 6'b111010;
		color_arr[3055] = 6'b111010;
		color_arr[3056] = 6'b111001;
		color_arr[3057] = 6'b000000;
		color_arr[3058] = 6'b000000;
		color_arr[3059] = 6'b000000;
		color_arr[3060] = 6'b000000;
		color_arr[3061] = 6'b000000;
		color_arr[3062] = 6'b000000;
		color_arr[3063] = 6'b000000;
		color_arr[3064] = 6'b000000;
		color_arr[3065] = 6'b000000;
		color_arr[3066] = 6'b000000;
		color_arr[3067] = 6'b000000;
		color_arr[3068] = 6'b000000;
		color_arr[3069] = 6'b000000;
		color_arr[3070] = 6'b000000;
		color_arr[3071] = 6'b000000;
		color_arr[3072] = 6'b000000;
		color_arr[3073] = 6'b000000;
		color_arr[3074] = 6'b000000;
		color_arr[3075] = 6'b000000;
		color_arr[3076] = 6'b000000;
		color_arr[3077] = 6'b000000;
		color_arr[3078] = 6'b000000;
		color_arr[3079] = 6'b000000;
		color_arr[3080] = 6'b000000;
		color_arr[3081] = 6'b000000;
		color_arr[3082] = 6'b000000;
		color_arr[3083] = 6'b000000;
		color_arr[3084] = 6'b000000;
		color_arr[3085] = 6'b000000;
		color_arr[3086] = 6'b000000;
		color_arr[3087] = 6'b111001;
		color_arr[3088] = 6'b111001;
		color_arr[3089] = 6'b111001;
		color_arr[3090] = 6'b111010;
		color_arr[3091] = 6'b111010;
		color_arr[3092] = 6'b111010;
		color_arr[3093] = 6'b111010;
		color_arr[3094] = 6'b111010;
		color_arr[3095] = 6'b111010;
		color_arr[3096] = 6'b111010;
		color_arr[3097] = 6'b111010;
		color_arr[3098] = 6'b111010;
		color_arr[3099] = 6'b111001;
		color_arr[3100] = 6'b111110;
		color_arr[3101] = 6'b111110;
		color_arr[3102] = 6'b111110;
		color_arr[3103] = 6'b111010;
		color_arr[3104] = 6'b111010;
		color_arr[3105] = 6'b111001;
		color_arr[3106] = 6'b111001;
		color_arr[3107] = 6'b111001;
		color_arr[3108] = 6'b111001;
		color_arr[3109] = 6'b111110;
		color_arr[3110] = 6'b111110;
		color_arr[3111] = 6'b111110;
		color_arr[3112] = 6'b111110;
		color_arr[3113] = 6'b111110;
		color_arr[3114] = 6'b111110;
		color_arr[3115] = 6'b111010;
		color_arr[3116] = 6'b111010;
		color_arr[3117] = 6'b111010;
		color_arr[3118] = 6'b111010;
		color_arr[3119] = 6'b111010;
		color_arr[3120] = 6'b111001;
		color_arr[3121] = 6'b000000;
		color_arr[3122] = 6'b000000;
		color_arr[3123] = 6'b000000;
		color_arr[3124] = 6'b000000;
		color_arr[3125] = 6'b000000;
		color_arr[3126] = 6'b000000;
		color_arr[3127] = 6'b000000;
		color_arr[3128] = 6'b000000;
		color_arr[3129] = 6'b000000;
		color_arr[3130] = 6'b000000;
		color_arr[3131] = 6'b000000;
		color_arr[3132] = 6'b000000;
		color_arr[3133] = 6'b000000;
		color_arr[3134] = 6'b000000;
		color_arr[3135] = 6'b000000;
		color_arr[3136] = 6'b000000;
		color_arr[3137] = 6'b000000;
		color_arr[3138] = 6'b000000;
		color_arr[3139] = 6'b000000;
		color_arr[3140] = 6'b000000;
		color_arr[3141] = 6'b000000;
		color_arr[3142] = 6'b000000;
		color_arr[3143] = 6'b000000;
		color_arr[3144] = 6'b000000;
		color_arr[3145] = 6'b000000;
		color_arr[3146] = 6'b000000;
		color_arr[3147] = 6'b000000;
		color_arr[3148] = 6'b000000;
		color_arr[3149] = 6'b000000;
		color_arr[3150] = 6'b000000;
		color_arr[3151] = 6'b111001;
		color_arr[3152] = 6'b111001;
		color_arr[3153] = 6'b111001;
		color_arr[3154] = 6'b111001;
		color_arr[3155] = 6'b111001;
		color_arr[3156] = 6'b111010;
		color_arr[3157] = 6'b111010;
		color_arr[3158] = 6'b111010;
		color_arr[3159] = 6'b111010;
		color_arr[3160] = 6'b111010;
		color_arr[3161] = 6'b111010;
		color_arr[3162] = 6'b111111;
		color_arr[3163] = 6'b111110;
		color_arr[3164] = 6'b111110;
		color_arr[3165] = 6'b111110;
		color_arr[3166] = 6'b111110;
		color_arr[3167] = 6'b111110;
		color_arr[3168] = 6'b111010;
		color_arr[3169] = 6'b111010;
		color_arr[3170] = 6'b111001;
		color_arr[3171] = 6'b111001;
		color_arr[3172] = 6'b111001;
		color_arr[3173] = 6'b111001;
		color_arr[3174] = 6'b111001;
		color_arr[3175] = 6'b111001;
		color_arr[3176] = 6'b111010;
		color_arr[3177] = 6'b111010;
		color_arr[3178] = 6'b111010;
		color_arr[3179] = 6'b111010;
		color_arr[3180] = 6'b111010;
		color_arr[3181] = 6'b111010;
		color_arr[3182] = 6'b111010;
		color_arr[3183] = 6'b111001;
		color_arr[3184] = 6'b111001;
		color_arr[3185] = 6'b000000;
		color_arr[3186] = 6'b000000;
		color_arr[3187] = 6'b000000;
		color_arr[3188] = 6'b000000;
		color_arr[3189] = 6'b000000;
		color_arr[3190] = 6'b000000;
		color_arr[3191] = 6'b000000;
		color_arr[3192] = 6'b000000;
		color_arr[3193] = 6'b000000;
		color_arr[3194] = 6'b000000;
		color_arr[3195] = 6'b000000;
		color_arr[3196] = 6'b000000;
		color_arr[3197] = 6'b000000;
		color_arr[3198] = 6'b000000;
		color_arr[3199] = 6'b000000;
		color_arr[3200] = 6'b000000;
		color_arr[3201] = 6'b000000;
		color_arr[3202] = 6'b000000;
		color_arr[3203] = 6'b000000;
		color_arr[3204] = 6'b000000;
		color_arr[3205] = 6'b000000;
		color_arr[3206] = 6'b000000;
		color_arr[3207] = 6'b000000;
		color_arr[3208] = 6'b000000;
		color_arr[3209] = 6'b000000;
		color_arr[3210] = 6'b000000;
		color_arr[3211] = 6'b000000;
		color_arr[3212] = 6'b000000;
		color_arr[3213] = 6'b000000;
		color_arr[3214] = 6'b000000;
		color_arr[3215] = 6'b000000;
		color_arr[3216] = 6'b111001;
		color_arr[3217] = 6'b111001;
		color_arr[3218] = 6'b111001;
		color_arr[3219] = 6'b111001;
		color_arr[3220] = 6'b111001;
		color_arr[3221] = 6'b111001;
		color_arr[3222] = 6'b111010;
		color_arr[3223] = 6'b111010;
		color_arr[3224] = 6'b111010;
		color_arr[3225] = 6'b111111;
		color_arr[3226] = 6'b111111;
		color_arr[3227] = 6'b111110;
		color_arr[3228] = 6'b111110;
		color_arr[3229] = 6'b111110;
		color_arr[3230] = 6'b111110;
		color_arr[3231] = 6'b111110;
		color_arr[3232] = 6'b111110;
		color_arr[3233] = 6'b111010;
		color_arr[3234] = 6'b111010;
		color_arr[3235] = 6'b111001;
		color_arr[3236] = 6'b111001;
		color_arr[3237] = 6'b111001;
		color_arr[3238] = 6'b111001;
		color_arr[3239] = 6'b111001;
		color_arr[3240] = 6'b111001;
		color_arr[3241] = 6'b111001;
		color_arr[3242] = 6'b111001;
		color_arr[3243] = 6'b111001;
		color_arr[3244] = 6'b111001;
		color_arr[3245] = 6'b111001;
		color_arr[3246] = 6'b111001;
		color_arr[3247] = 6'b111001;
		color_arr[3248] = 6'b111001;
		color_arr[3249] = 6'b000000;
		color_arr[3250] = 6'b000000;
		color_arr[3251] = 6'b000000;
		color_arr[3252] = 6'b000000;
		color_arr[3253] = 6'b000000;
		color_arr[3254] = 6'b000000;
		color_arr[3255] = 6'b000000;
		color_arr[3256] = 6'b000000;
		color_arr[3257] = 6'b000000;
		color_arr[3258] = 6'b000000;
		color_arr[3259] = 6'b000000;
		color_arr[3260] = 6'b000000;
		color_arr[3261] = 6'b000000;
		color_arr[3262] = 6'b000000;
		color_arr[3263] = 6'b000000;
		color_arr[3264] = 6'b000000;
		color_arr[3265] = 6'b000000;
		color_arr[3266] = 6'b000000;
		color_arr[3267] = 6'b000000;
		color_arr[3268] = 6'b000000;
		color_arr[3269] = 6'b000000;
		color_arr[3270] = 6'b000000;
		color_arr[3271] = 6'b000000;
		color_arr[3272] = 6'b000000;
		color_arr[3273] = 6'b000000;
		color_arr[3274] = 6'b000000;
		color_arr[3275] = 6'b000000;
		color_arr[3276] = 6'b000000;
		color_arr[3277] = 6'b000000;
		color_arr[3278] = 6'b000000;
		color_arr[3279] = 6'b000000;
		color_arr[3280] = 6'b000000;
		color_arr[3281] = 6'b000000;
		color_arr[3282] = 6'b111001;
		color_arr[3283] = 6'b111001;
		color_arr[3284] = 6'b111001;
		color_arr[3285] = 6'b111001;
		color_arr[3286] = 6'b111001;
		color_arr[3287] = 6'b111010;
		color_arr[3288] = 6'b111111;
		color_arr[3289] = 6'b111111;
		color_arr[3290] = 6'b111111;
		color_arr[3291] = 6'b111111;
		color_arr[3292] = 6'b111111;
		color_arr[3293] = 6'b111110;
		color_arr[3294] = 6'b111110;
		color_arr[3295] = 6'b111110;
		color_arr[3296] = 6'b111110;
		color_arr[3297] = 6'b111110;
		color_arr[3298] = 6'b111010;
		color_arr[3299] = 6'b111010;
		color_arr[3300] = 6'b111001;
		color_arr[3301] = 6'b111001;
		color_arr[3302] = 6'b111001;
		color_arr[3303] = 6'b111001;
		color_arr[3304] = 6'b111001;
		color_arr[3305] = 6'b111001;
		color_arr[3306] = 6'b111001;
		color_arr[3307] = 6'b111001;
		color_arr[3308] = 6'b111001;
		color_arr[3309] = 6'b111001;
		color_arr[3310] = 6'b111001;
		color_arr[3311] = 6'b111001;
		color_arr[3312] = 6'b111001;
		color_arr[3313] = 6'b000000;
		color_arr[3314] = 6'b000000;
		color_arr[3315] = 6'b000000;
		color_arr[3316] = 6'b000000;
		color_arr[3317] = 6'b000000;
		color_arr[3318] = 6'b000000;
		color_arr[3319] = 6'b000000;
		color_arr[3320] = 6'b000000;
		color_arr[3321] = 6'b000000;
		color_arr[3322] = 6'b000000;
		color_arr[3323] = 6'b000000;
		color_arr[3324] = 6'b000000;
		color_arr[3325] = 6'b000000;
		color_arr[3326] = 6'b000000;
		color_arr[3327] = 6'b000000;
		color_arr[3328] = 6'b000000;
		color_arr[3329] = 6'b000000;
		color_arr[3330] = 6'b000000;
		color_arr[3331] = 6'b000000;
		color_arr[3332] = 6'b000000;
		color_arr[3333] = 6'b000000;
		color_arr[3334] = 6'b000000;
		color_arr[3335] = 6'b000000;
		color_arr[3336] = 6'b000000;
		color_arr[3337] = 6'b000000;
		color_arr[3338] = 6'b000000;
		color_arr[3339] = 6'b000000;
		color_arr[3340] = 6'b000000;
		color_arr[3341] = 6'b000000;
		color_arr[3342] = 6'b000000;
		color_arr[3343] = 6'b000000;
		color_arr[3344] = 6'b000000;
		color_arr[3345] = 6'b000000;
		color_arr[3346] = 6'b000000;
		color_arr[3347] = 6'b000000;
		color_arr[3348] = 6'b000000;
		color_arr[3349] = 6'b111001;
		color_arr[3350] = 6'b111001;
		color_arr[3351] = 6'b111001;
		color_arr[3352] = 6'b111110;
		color_arr[3353] = 6'b111111;
		color_arr[3354] = 6'b111111;
		color_arr[3355] = 6'b111111;
		color_arr[3356] = 6'b111111;
		color_arr[3357] = 6'b111111;
		color_arr[3358] = 6'b111111;
		color_arr[3359] = 6'b111110;
		color_arr[3360] = 6'b111110;
		color_arr[3361] = 6'b111110;
		color_arr[3362] = 6'b111010;
		color_arr[3363] = 6'b111010;
		color_arr[3364] = 6'b111001;
		color_arr[3365] = 6'b111001;
		color_arr[3366] = 6'b111001;
		color_arr[3367] = 6'b111001;
		color_arr[3368] = 6'b111010;
		color_arr[3369] = 6'b111010;
		color_arr[3370] = 6'b111010;
		color_arr[3371] = 6'b111010;
		color_arr[3372] = 6'b111001;
		color_arr[3373] = 6'b111001;
		color_arr[3374] = 6'b111001;
		color_arr[3375] = 6'b111001;
		color_arr[3376] = 6'b000000;
		color_arr[3377] = 6'b000000;
		color_arr[3378] = 6'b000000;
		color_arr[3379] = 6'b000000;
		color_arr[3380] = 6'b000000;
		color_arr[3381] = 6'b000000;
		color_arr[3382] = 6'b000000;
		color_arr[3383] = 6'b000000;
		color_arr[3384] = 6'b000000;
		color_arr[3385] = 6'b000000;
		color_arr[3386] = 6'b000000;
		color_arr[3387] = 6'b000000;
		color_arr[3388] = 6'b000000;
		color_arr[3389] = 6'b000000;
		color_arr[3390] = 6'b000000;
		color_arr[3391] = 6'b000000;
		color_arr[3392] = 6'b000000;
		color_arr[3393] = 6'b000000;
		color_arr[3394] = 6'b000000;
		color_arr[3395] = 6'b000000;
		color_arr[3396] = 6'b000000;
		color_arr[3397] = 6'b000000;
		color_arr[3398] = 6'b000000;
		color_arr[3399] = 6'b000000;
		color_arr[3400] = 6'b000000;
		color_arr[3401] = 6'b000000;
		color_arr[3402] = 6'b000000;
		color_arr[3403] = 6'b000000;
		color_arr[3404] = 6'b000000;
		color_arr[3405] = 6'b000000;
		color_arr[3406] = 6'b000000;
		color_arr[3407] = 6'b000000;
		color_arr[3408] = 6'b000000;
		color_arr[3409] = 6'b000000;
		color_arr[3410] = 6'b000000;
		color_arr[3411] = 6'b000000;
		color_arr[3412] = 6'b000000;
		color_arr[3413] = 6'b000000;
		color_arr[3414] = 6'b000000;
		color_arr[3415] = 6'b111001;
		color_arr[3416] = 6'b111111;
		color_arr[3417] = 6'b111110;
		color_arr[3418] = 6'b111111;
		color_arr[3419] = 6'b111110;
		color_arr[3420] = 6'b111110;
		color_arr[3421] = 6'b111111;
		color_arr[3422] = 6'b111111;
		color_arr[3423] = 6'b111111;
		color_arr[3424] = 6'b111110;
		color_arr[3425] = 6'b111110;
		color_arr[3426] = 6'b111010;
		color_arr[3427] = 6'b111001;
		color_arr[3428] = 6'b111001;
		color_arr[3429] = 6'b111010;
		color_arr[3430] = 6'b111010;
		color_arr[3431] = 6'b111010;
		color_arr[3432] = 6'b111010;
		color_arr[3433] = 6'b111010;
		color_arr[3434] = 6'b111010;
		color_arr[3435] = 6'b111010;
		color_arr[3436] = 6'b111010;
		color_arr[3437] = 6'b111001;
		color_arr[3438] = 6'b111001;
		color_arr[3439] = 6'b111001;
		color_arr[3440] = 6'b000000;
		color_arr[3441] = 6'b000000;
		color_arr[3442] = 6'b000000;
		color_arr[3443] = 6'b000000;
		color_arr[3444] = 6'b000000;
		color_arr[3445] = 6'b000000;
		color_arr[3446] = 6'b000000;
		color_arr[3447] = 6'b000000;
		color_arr[3448] = 6'b000000;
		color_arr[3449] = 6'b000000;
		color_arr[3450] = 6'b000000;
		color_arr[3451] = 6'b000000;
		color_arr[3452] = 6'b000000;
		color_arr[3453] = 6'b000000;
		color_arr[3454] = 6'b000000;
		color_arr[3455] = 6'b000000;
		color_arr[3456] = 6'b000000;
		color_arr[3457] = 6'b000000;
		color_arr[3458] = 6'b000000;
		color_arr[3459] = 6'b000000;
		color_arr[3460] = 6'b000000;
		color_arr[3461] = 6'b000000;
		color_arr[3462] = 6'b000000;
		color_arr[3463] = 6'b000000;
		color_arr[3464] = 6'b000000;
		color_arr[3465] = 6'b000000;
		color_arr[3466] = 6'b000000;
		color_arr[3467] = 6'b000000;
		color_arr[3468] = 6'b000000;
		color_arr[3469] = 6'b000000;
		color_arr[3470] = 6'b000000;
		color_arr[3471] = 6'b000000;
		color_arr[3472] = 6'b000000;
		color_arr[3473] = 6'b000000;
		color_arr[3474] = 6'b000000;
		color_arr[3475] = 6'b000000;
		color_arr[3476] = 6'b000000;
		color_arr[3477] = 6'b000000;
		color_arr[3478] = 6'b000000;
		color_arr[3479] = 6'b000000;
		color_arr[3480] = 6'b010101;
		color_arr[3481] = 6'b111111;
		color_arr[3482] = 6'b111110;
		color_arr[3483] = 6'b111111;
		color_arr[3484] = 6'b111110;
		color_arr[3485] = 6'b111111;
		color_arr[3486] = 6'b111111;
		color_arr[3487] = 6'b111010;
		color_arr[3488] = 6'b111010;
		color_arr[3489] = 6'b111010;
		color_arr[3490] = 6'b111001;
		color_arr[3491] = 6'b111001;
		color_arr[3492] = 6'b111001;
		color_arr[3493] = 6'b111001;
		color_arr[3494] = 6'b111010;
		color_arr[3495] = 6'b111010;
		color_arr[3496] = 6'b111010;
		color_arr[3497] = 6'b111010;
		color_arr[3498] = 6'b111010;
		color_arr[3499] = 6'b111010;
		color_arr[3500] = 6'b111001;
		color_arr[3501] = 6'b111001;
		color_arr[3502] = 6'b111001;
		color_arr[3503] = 6'b111001;
		color_arr[3504] = 6'b000000;
		color_arr[3505] = 6'b000000;
		color_arr[3506] = 6'b000000;
		color_arr[3507] = 6'b000000;
		color_arr[3508] = 6'b000000;
		color_arr[3509] = 6'b000000;
		color_arr[3510] = 6'b000000;
		color_arr[3511] = 6'b000000;
		color_arr[3512] = 6'b000000;
		color_arr[3513] = 6'b000000;
		color_arr[3514] = 6'b000000;
		color_arr[3515] = 6'b000000;
		color_arr[3516] = 6'b000000;
		color_arr[3517] = 6'b000000;
		color_arr[3518] = 6'b000000;
		color_arr[3519] = 6'b000000;
		color_arr[3520] = 6'b000000;
		color_arr[3521] = 6'b000000;
		color_arr[3522] = 6'b000000;
		color_arr[3523] = 6'b000000;
		color_arr[3524] = 6'b000000;
		color_arr[3525] = 6'b000000;
		color_arr[3526] = 6'b000000;
		color_arr[3527] = 6'b000000;
		color_arr[3528] = 6'b000000;
		color_arr[3529] = 6'b000000;
		color_arr[3530] = 6'b000000;
		color_arr[3531] = 6'b000000;
		color_arr[3532] = 6'b000000;
		color_arr[3533] = 6'b000000;
		color_arr[3534] = 6'b000000;
		color_arr[3535] = 6'b000000;
		color_arr[3536] = 6'b000000;
		color_arr[3537] = 6'b000000;
		color_arr[3538] = 6'b000000;
		color_arr[3539] = 6'b000000;
		color_arr[3540] = 6'b000000;
		color_arr[3541] = 6'b000000;
		color_arr[3542] = 6'b000000;
		color_arr[3543] = 6'b000000;
		color_arr[3544] = 6'b000000;
		color_arr[3545] = 6'b010101;
		color_arr[3546] = 6'b111110;
		color_arr[3547] = 6'b010101;
		color_arr[3548] = 6'b111110;
		color_arr[3549] = 6'b010101;
		color_arr[3550] = 6'b111010;
		color_arr[3551] = 6'b111010;
		color_arr[3552] = 6'b111010;
		color_arr[3553] = 6'b111010;
		color_arr[3554] = 6'b111010;
		color_arr[3555] = 6'b111001;
		color_arr[3556] = 6'b111001;
		color_arr[3557] = 6'b111001;
		color_arr[3558] = 6'b111001;
		color_arr[3559] = 6'b111001;
		color_arr[3560] = 6'b111001;
		color_arr[3561] = 6'b111001;
		color_arr[3562] = 6'b111001;
		color_arr[3563] = 6'b111001;
		color_arr[3564] = 6'b111001;
		color_arr[3565] = 6'b111001;
		color_arr[3566] = 6'b111001;
		color_arr[3567] = 6'b000000;
		color_arr[3568] = 6'b000000;
		color_arr[3569] = 6'b000000;
		color_arr[3570] = 6'b000000;
		color_arr[3571] = 6'b000000;
		color_arr[3572] = 6'b000000;
		color_arr[3573] = 6'b000000;
		color_arr[3574] = 6'b000000;
		color_arr[3575] = 6'b000000;
		color_arr[3576] = 6'b000000;
		color_arr[3577] = 6'b000000;
		color_arr[3578] = 6'b000000;
		color_arr[3579] = 6'b000000;
		color_arr[3580] = 6'b000000;
		color_arr[3581] = 6'b000000;
		color_arr[3582] = 6'b000000;
		color_arr[3583] = 6'b000000;
		color_arr[3584] = 6'b000000;
		color_arr[3585] = 6'b000000;
		color_arr[3586] = 6'b000000;
		color_arr[3587] = 6'b000000;
		color_arr[3588] = 6'b000000;
		color_arr[3589] = 6'b000000;
		color_arr[3590] = 6'b000000;
		color_arr[3591] = 6'b000000;
		color_arr[3592] = 6'b000000;
		color_arr[3593] = 6'b000000;
		color_arr[3594] = 6'b000000;
		color_arr[3595] = 6'b000000;
		color_arr[3596] = 6'b000000;
		color_arr[3597] = 6'b000000;
		color_arr[3598] = 6'b000000;
		color_arr[3599] = 6'b000000;
		color_arr[3600] = 6'b000000;
		color_arr[3601] = 6'b000000;
		color_arr[3602] = 6'b000000;
		color_arr[3603] = 6'b000000;
		color_arr[3604] = 6'b000000;
		color_arr[3605] = 6'b000000;
		color_arr[3606] = 6'b000000;
		color_arr[3607] = 6'b000000;
		color_arr[3608] = 6'b000000;
		color_arr[3609] = 6'b000000;
		color_arr[3610] = 6'b000000;
		color_arr[3611] = 6'b111010;
		color_arr[3612] = 6'b111010;
		color_arr[3613] = 6'b111010;
		color_arr[3614] = 6'b111010;
		color_arr[3615] = 6'b111010;
		color_arr[3616] = 6'b111010;
		color_arr[3617] = 6'b111010;
		color_arr[3618] = 6'b111010;
		color_arr[3619] = 6'b000000;
		color_arr[3620] = 6'b111001;
		color_arr[3621] = 6'b111001;
		color_arr[3622] = 6'b111001;
		color_arr[3623] = 6'b111001;
		color_arr[3624] = 6'b111001;
		color_arr[3625] = 6'b111001;
		color_arr[3626] = 6'b111001;
		color_arr[3627] = 6'b111001;
		color_arr[3628] = 6'b111001;
		color_arr[3629] = 6'b111001;
		color_arr[3630] = 6'b000000;
		color_arr[3631] = 6'b000000;
		color_arr[3632] = 6'b000000;
		color_arr[3633] = 6'b000000;
		color_arr[3634] = 6'b000000;
		color_arr[3635] = 6'b000000;
		color_arr[3636] = 6'b000000;
		color_arr[3637] = 6'b000000;
		color_arr[3638] = 6'b000000;
		color_arr[3639] = 6'b000000;
		color_arr[3640] = 6'b000000;
		color_arr[3641] = 6'b000000;
		color_arr[3642] = 6'b000000;
		color_arr[3643] = 6'b000000;
		color_arr[3644] = 6'b000000;
		color_arr[3645] = 6'b000000;
		color_arr[3646] = 6'b000000;
		color_arr[3647] = 6'b000000;
		color_arr[3648] = 6'b000000;
		color_arr[3649] = 6'b000000;
		color_arr[3650] = 6'b000000;
		color_arr[3651] = 6'b000000;
		color_arr[3652] = 6'b000000;
		color_arr[3653] = 6'b000000;
		color_arr[3654] = 6'b000000;
		color_arr[3655] = 6'b000000;
		color_arr[3656] = 6'b000000;
		color_arr[3657] = 6'b000000;
		color_arr[3658] = 6'b000000;
		color_arr[3659] = 6'b000000;
		color_arr[3660] = 6'b000000;
		color_arr[3661] = 6'b000000;
		color_arr[3662] = 6'b000000;
		color_arr[3663] = 6'b000000;
		color_arr[3664] = 6'b000000;
		color_arr[3665] = 6'b000000;
		color_arr[3666] = 6'b000000;
		color_arr[3667] = 6'b000000;
		color_arr[3668] = 6'b000000;
		color_arr[3669] = 6'b000000;
		color_arr[3670] = 6'b000000;
		color_arr[3671] = 6'b000000;
		color_arr[3672] = 6'b000000;
		color_arr[3673] = 6'b000000;
		color_arr[3674] = 6'b000000;
		color_arr[3675] = 6'b000000;
		color_arr[3676] = 6'b111010;
		color_arr[3677] = 6'b111010;
		color_arr[3678] = 6'b111010;
		color_arr[3679] = 6'b111010;
		color_arr[3680] = 6'b111010;
		color_arr[3681] = 6'b010101;
		color_arr[3682] = 6'b000000;
		color_arr[3683] = 6'b000000;
		color_arr[3684] = 6'b000000;
		color_arr[3685] = 6'b000000;
		color_arr[3686] = 6'b000000;
		color_arr[3687] = 6'b111001;
		color_arr[3688] = 6'b111001;
		color_arr[3689] = 6'b111001;
		color_arr[3690] = 6'b111001;
		color_arr[3691] = 6'b111001;
		color_arr[3692] = 6'b111001;
		color_arr[3693] = 6'b000000;
		color_arr[3694] = 6'b000000;
		color_arr[3695] = 6'b000000;
		color_arr[3696] = 6'b000000;
		color_arr[3697] = 6'b000000;
		color_arr[3698] = 6'b000000;
		color_arr[3699] = 6'b000000;
		color_arr[3700] = 6'b000000;
		color_arr[3701] = 6'b000000;
		color_arr[3702] = 6'b000000;
		color_arr[3703] = 6'b000000;
		color_arr[3704] = 6'b000000;
		color_arr[3705] = 6'b000000;
		color_arr[3706] = 6'b000000;
		color_arr[3707] = 6'b000000;
		color_arr[3708] = 6'b000000;
		color_arr[3709] = 6'b000000;
		color_arr[3710] = 6'b000000;
		color_arr[3711] = 6'b000000;
		color_arr[3712] = 6'b000000;
		color_arr[3713] = 6'b000000;
		color_arr[3714] = 6'b000000;
		color_arr[3715] = 6'b000000;
		color_arr[3716] = 6'b000000;
		color_arr[3717] = 6'b000000;
		color_arr[3718] = 6'b000000;
		color_arr[3719] = 6'b000000;
		color_arr[3720] = 6'b000000;
		color_arr[3721] = 6'b000000;
		color_arr[3722] = 6'b000000;
		color_arr[3723] = 6'b000000;
		color_arr[3724] = 6'b000000;
		color_arr[3725] = 6'b000000;
		color_arr[3726] = 6'b000000;
		color_arr[3727] = 6'b000000;
		color_arr[3728] = 6'b000000;
		color_arr[3729] = 6'b000000;
		color_arr[3730] = 6'b000000;
		color_arr[3731] = 6'b000000;
		color_arr[3732] = 6'b000000;
		color_arr[3733] = 6'b000000;
		color_arr[3734] = 6'b000000;
		color_arr[3735] = 6'b000000;
		color_arr[3736] = 6'b000000;
		color_arr[3737] = 6'b000000;
		color_arr[3738] = 6'b000000;
		color_arr[3739] = 6'b000000;
		color_arr[3740] = 6'b000000;
		color_arr[3741] = 6'b000000;
		color_arr[3742] = 6'b111010;
		color_arr[3743] = 6'b010101;
		color_arr[3744] = 6'b000000;
		color_arr[3745] = 6'b000000;
		color_arr[3746] = 6'b000000;
		color_arr[3747] = 6'b000000;
		color_arr[3748] = 6'b000000;
		color_arr[3749] = 6'b000000;
		color_arr[3750] = 6'b000000;
		color_arr[3751] = 6'b000000;
		color_arr[3752] = 6'b000000;
		color_arr[3753] = 6'b000000;
		color_arr[3754] = 6'b000000;
		color_arr[3755] = 6'b000000;
		color_arr[3756] = 6'b000000;
		color_arr[3757] = 6'b000000;
		color_arr[3758] = 6'b000000;
		color_arr[3759] = 6'b000000;
		color_arr[3760] = 6'b000000;
		color_arr[3761] = 6'b000000;
		color_arr[3762] = 6'b000000;
		color_arr[3763] = 6'b000000;
		color_arr[3764] = 6'b000000;
		color_arr[3765] = 6'b000000;
		color_arr[3766] = 6'b000000;
		color_arr[3767] = 6'b000000;
		color_arr[3768] = 6'b000000;
		color_arr[3769] = 6'b000000;
		color_arr[3770] = 6'b000000;
		color_arr[3771] = 6'b000000;
		color_arr[3772] = 6'b000000;
		color_arr[3773] = 6'b000000;
		color_arr[3774] = 6'b000000;
		color_arr[3775] = 6'b000000;
		color_arr[3776] = 6'b000000;
		color_arr[3777] = 6'b000000;
		color_arr[3778] = 6'b000000;
		color_arr[3779] = 6'b000000;
		color_arr[3780] = 6'b000000;
		color_arr[3781] = 6'b000000;
		color_arr[3782] = 6'b000000;
		color_arr[3783] = 6'b000000;
		color_arr[3784] = 6'b000000;
		color_arr[3785] = 6'b000000;
		color_arr[3786] = 6'b000000;
		color_arr[3787] = 6'b000000;
		color_arr[3788] = 6'b000000;
		color_arr[3789] = 6'b000000;
		color_arr[3790] = 6'b000000;
		color_arr[3791] = 6'b000000;
		color_arr[3792] = 6'b000000;
		color_arr[3793] = 6'b000000;
		color_arr[3794] = 6'b000000;
		color_arr[3795] = 6'b000000;
		color_arr[3796] = 6'b000000;
		color_arr[3797] = 6'b000000;
		color_arr[3798] = 6'b000000;
		color_arr[3799] = 6'b000000;
		color_arr[3800] = 6'b000000;
		color_arr[3801] = 6'b000000;
		color_arr[3802] = 6'b000000;
		color_arr[3803] = 6'b000000;
		color_arr[3804] = 6'b000000;
		color_arr[3805] = 6'b000000;
		color_arr[3806] = 6'b000000;
		color_arr[3807] = 6'b000000;
		color_arr[3808] = 6'b000000;
		color_arr[3809] = 6'b000000;
		color_arr[3810] = 6'b000000;
		color_arr[3811] = 6'b000000;
		color_arr[3812] = 6'b000000;
		color_arr[3813] = 6'b000000;
		color_arr[3814] = 6'b000000;
		color_arr[3815] = 6'b000000;
		color_arr[3816] = 6'b000000;
		color_arr[3817] = 6'b000000;
		color_arr[3818] = 6'b000000;
		color_arr[3819] = 6'b000000;
		color_arr[3820] = 6'b000000;
		color_arr[3821] = 6'b000000;
		color_arr[3822] = 6'b000000;
		color_arr[3823] = 6'b000000;
		color_arr[3824] = 6'b000000;
		color_arr[3825] = 6'b000000;
		color_arr[3826] = 6'b000000;
		color_arr[3827] = 6'b000000;
		color_arr[3828] = 6'b000000;
		color_arr[3829] = 6'b000000;
		color_arr[3830] = 6'b000000;
		color_arr[3831] = 6'b000000;
		color_arr[3832] = 6'b000000;
		color_arr[3833] = 6'b000000;
		color_arr[3834] = 6'b000000;
		color_arr[3835] = 6'b000000;
		color_arr[3836] = 6'b000000;
		color_arr[3837] = 6'b000000;
		color_arr[3838] = 6'b000000;
		color_arr[3839] = 6'b000000;
		color_arr[3840] = 6'b000000;
		color_arr[3841] = 6'b000000;
		color_arr[3842] = 6'b000000;
		color_arr[3843] = 6'b000000;
		color_arr[3844] = 6'b000000;
		color_arr[3845] = 6'b000000;
		color_arr[3846] = 6'b000000;
		color_arr[3847] = 6'b000000;
		color_arr[3848] = 6'b000000;
		color_arr[3849] = 6'b000000;
		color_arr[3850] = 6'b000000;
		color_arr[3851] = 6'b000000;
		color_arr[3852] = 6'b000000;
		color_arr[3853] = 6'b000000;
		color_arr[3854] = 6'b000000;
		color_arr[3855] = 6'b000000;
		color_arr[3856] = 6'b000000;
		color_arr[3857] = 6'b000000;
		color_arr[3858] = 6'b000000;
		color_arr[3859] = 6'b000000;
		color_arr[3860] = 6'b000000;
		color_arr[3861] = 6'b000000;
		color_arr[3862] = 6'b000000;
		color_arr[3863] = 6'b000000;
		color_arr[3864] = 6'b000000;
		color_arr[3865] = 6'b000000;
		color_arr[3866] = 6'b000000;
		color_arr[3867] = 6'b000000;
		color_arr[3868] = 6'b000000;
		color_arr[3869] = 6'b000000;
		color_arr[3870] = 6'b000000;
		color_arr[3871] = 6'b000000;
		color_arr[3872] = 6'b000000;
		color_arr[3873] = 6'b000000;
		color_arr[3874] = 6'b000000;
		color_arr[3875] = 6'b000000;
		color_arr[3876] = 6'b000000;
		color_arr[3877] = 6'b000000;
		color_arr[3878] = 6'b000000;
		color_arr[3879] = 6'b000000;
		color_arr[3880] = 6'b000000;
		color_arr[3881] = 6'b000000;
		color_arr[3882] = 6'b000000;
		color_arr[3883] = 6'b000000;
		color_arr[3884] = 6'b000000;
		color_arr[3885] = 6'b000000;
		color_arr[3886] = 6'b000000;
		color_arr[3887] = 6'b000000;
		color_arr[3888] = 6'b000000;
		color_arr[3889] = 6'b000000;
		color_arr[3890] = 6'b000000;
		color_arr[3891] = 6'b000000;
		color_arr[3892] = 6'b000000;
		color_arr[3893] = 6'b000000;
		color_arr[3894] = 6'b000000;
		color_arr[3895] = 6'b000000;
		color_arr[3896] = 6'b000000;
		color_arr[3897] = 6'b000000;
		color_arr[3898] = 6'b000000;
		color_arr[3899] = 6'b000000;
		color_arr[3900] = 6'b000000;
		color_arr[3901] = 6'b000000;
		color_arr[3902] = 6'b000000;
		color_arr[3903] = 6'b000000;
		color_arr[3904] = 6'b000000;
		color_arr[3905] = 6'b000000;
		color_arr[3906] = 6'b000000;
		color_arr[3907] = 6'b000000;
		color_arr[3908] = 6'b000000;
		color_arr[3909] = 6'b000000;
		color_arr[3910] = 6'b000000;
		color_arr[3911] = 6'b000000;
		color_arr[3912] = 6'b000000;
		color_arr[3913] = 6'b000000;
		color_arr[3914] = 6'b000000;
		color_arr[3915] = 6'b000000;
		color_arr[3916] = 6'b000000;
		color_arr[3917] = 6'b000000;
		color_arr[3918] = 6'b000000;
		color_arr[3919] = 6'b000000;
		color_arr[3920] = 6'b000000;
		color_arr[3921] = 6'b000000;
		color_arr[3922] = 6'b000000;
		color_arr[3923] = 6'b000000;
		color_arr[3924] = 6'b000000;
		color_arr[3925] = 6'b000000;
		color_arr[3926] = 6'b000000;
		color_arr[3927] = 6'b000000;
		color_arr[3928] = 6'b000000;
		color_arr[3929] = 6'b000000;
		color_arr[3930] = 6'b000000;
		color_arr[3931] = 6'b000000;
		color_arr[3932] = 6'b000000;
		color_arr[3933] = 6'b000000;
		color_arr[3934] = 6'b000000;
		color_arr[3935] = 6'b000000;
		color_arr[3936] = 6'b000000;
		color_arr[3937] = 6'b000000;
		color_arr[3938] = 6'b000000;
		color_arr[3939] = 6'b000000;
		color_arr[3940] = 6'b000000;
		color_arr[3941] = 6'b000000;
		color_arr[3942] = 6'b000000;
		color_arr[3943] = 6'b000000;
		color_arr[3944] = 6'b000000;
		color_arr[3945] = 6'b000000;
		color_arr[3946] = 6'b000000;
		color_arr[3947] = 6'b000000;
		color_arr[3948] = 6'b000000;
		color_arr[3949] = 6'b000000;
		color_arr[3950] = 6'b000000;
		color_arr[3951] = 6'b000000;
		color_arr[3952] = 6'b000000;
		color_arr[3953] = 6'b000000;
		color_arr[3954] = 6'b000000;
		color_arr[3955] = 6'b000000;
		color_arr[3956] = 6'b000000;
		color_arr[3957] = 6'b000000;
		color_arr[3958] = 6'b000000;
		color_arr[3959] = 6'b000000;
		color_arr[3960] = 6'b000000;
		color_arr[3961] = 6'b000000;
		color_arr[3962] = 6'b000000;
		color_arr[3963] = 6'b000000;
		color_arr[3964] = 6'b000000;
		color_arr[3965] = 6'b000000;
		color_arr[3966] = 6'b000000;
		color_arr[3967] = 6'b000000;
		color_arr[3968] = 6'b000000;
		color_arr[3969] = 6'b000000;
		color_arr[3970] = 6'b000000;
		color_arr[3971] = 6'b000000;
		color_arr[3972] = 6'b000000;
		color_arr[3973] = 6'b000000;
		color_arr[3974] = 6'b000000;
		color_arr[3975] = 6'b000000;
		color_arr[3976] = 6'b000000;
		color_arr[3977] = 6'b000000;
		color_arr[3978] = 6'b000000;
		color_arr[3979] = 6'b000000;
		color_arr[3980] = 6'b000000;
		color_arr[3981] = 6'b000000;
		color_arr[3982] = 6'b000000;
		color_arr[3983] = 6'b000000;
		color_arr[3984] = 6'b000000;
		color_arr[3985] = 6'b000000;
		color_arr[3986] = 6'b000000;
		color_arr[3987] = 6'b000000;
		color_arr[3988] = 6'b000000;
		color_arr[3989] = 6'b000000;
		color_arr[3990] = 6'b000000;
		color_arr[3991] = 6'b000000;
		color_arr[3992] = 6'b000000;
		color_arr[3993] = 6'b000000;
		color_arr[3994] = 6'b000000;
		color_arr[3995] = 6'b000000;
		color_arr[3996] = 6'b000000;
		color_arr[3997] = 6'b000000;
		color_arr[3998] = 6'b000000;
		color_arr[3999] = 6'b000000;
		color_arr[4000] = 6'b000000;
		color_arr[4001] = 6'b000000;
		color_arr[4002] = 6'b000000;
		color_arr[4003] = 6'b000000;
		color_arr[4004] = 6'b000000;
		color_arr[4005] = 6'b000000;
		color_arr[4006] = 6'b000000;
		color_arr[4007] = 6'b000000;
		color_arr[4008] = 6'b000000;
		color_arr[4009] = 6'b000000;
		color_arr[4010] = 6'b000000;
		color_arr[4011] = 6'b000000;
		color_arr[4012] = 6'b000000;
		color_arr[4013] = 6'b000000;
		color_arr[4014] = 6'b000000;
		color_arr[4015] = 6'b000000;
		color_arr[4016] = 6'b000000;
		color_arr[4017] = 6'b000000;
		color_arr[4018] = 6'b000000;
		color_arr[4019] = 6'b000000;
		color_arr[4020] = 6'b000000;
		color_arr[4021] = 6'b000000;
		color_arr[4022] = 6'b000000;
		color_arr[4023] = 6'b000000;
		color_arr[4024] = 6'b000000;
		color_arr[4025] = 6'b000000;
		color_arr[4026] = 6'b000000;
		color_arr[4027] = 6'b000000;
		color_arr[4028] = 6'b000000;
		color_arr[4029] = 6'b000000;
		color_arr[4030] = 6'b000000;
		color_arr[4031] = 6'b000000;
		color_arr[4032] = 6'b000000;
		color_arr[4033] = 6'b000000;
		color_arr[4034] = 6'b000000;
		color_arr[4035] = 6'b000000;
		color_arr[4036] = 6'b000000;
		color_arr[4037] = 6'b000000;
		color_arr[4038] = 6'b000000;
		color_arr[4039] = 6'b000000;
		color_arr[4040] = 6'b000000;
		color_arr[4041] = 6'b000000;
		color_arr[4042] = 6'b000000;
		color_arr[4043] = 6'b000000;
		color_arr[4044] = 6'b000000;
		color_arr[4045] = 6'b000000;
		color_arr[4046] = 6'b000000;
		color_arr[4047] = 6'b000000;
		color_arr[4048] = 6'b000000;
		color_arr[4049] = 6'b000000;
		color_arr[4050] = 6'b000000;
		color_arr[4051] = 6'b000000;
		color_arr[4052] = 6'b000000;
		color_arr[4053] = 6'b000000;
		color_arr[4054] = 6'b000000;
		color_arr[4055] = 6'b000000;
		color_arr[4056] = 6'b000000;
		color_arr[4057] = 6'b000000;
		color_arr[4058] = 6'b000000;
		color_arr[4059] = 6'b000000;
		color_arr[4060] = 6'b000000;
		color_arr[4061] = 6'b000000;
		color_arr[4062] = 6'b000000;
		color_arr[4063] = 6'b000000;
		color_arr[4064] = 6'b000000;
		color_arr[4065] = 6'b000000;
		color_arr[4066] = 6'b000000;
		color_arr[4067] = 6'b000000;
		color_arr[4068] = 6'b000000;
		color_arr[4069] = 6'b000000;
		color_arr[4070] = 6'b000000;
		color_arr[4071] = 6'b000000;
		color_arr[4072] = 6'b000000;
		color_arr[4073] = 6'b000000;
		color_arr[4074] = 6'b000000;
		color_arr[4075] = 6'b000000;
		color_arr[4076] = 6'b000000;
		color_arr[4077] = 6'b000000;
		color_arr[4078] = 6'b000000;
		color_arr[4079] = 6'b000000;
		color_arr[4080] = 6'b000000;
		color_arr[4081] = 6'b000000;
		color_arr[4082] = 6'b000000;
		color_arr[4083] = 6'b000000;
		color_arr[4084] = 6'b000000;
		color_arr[4085] = 6'b000000;
		color_arr[4086] = 6'b000000;
		color_arr[4087] = 6'b000000;
		color_arr[4088] = 6'b000000;
		color_arr[4089] = 6'b000000;
		color_arr[4090] = 6'b000000;
		color_arr[4091] = 6'b000000;
		color_arr[4092] = 6'b000000;
		color_arr[4093] = 6'b000000;
		color_arr[4094] = 6'b000000;
		color_arr[4095] = 6'b000000;
	end

	always @(posedge clk) begin
		color_out <= color_arr[addr];
	end
endmodule
