module sprite_rom (
	input clk,
	input [10:0] addr,
	output reg [5:0] color_out
);
	reg [7:0] color_arr [2047:0];

	initial begin
		color_arr[0] = 8'h0F;
		color_arr[1] = 8'h0F;
		color_arr[2] = 8'h0F;
		color_arr[3] = 8'h0F;
		color_arr[4] = 8'h0F;
		color_arr[5] = 8'h0F;
		color_arr[6] = 8'h0F;
		color_arr[7] = 8'h0F;
		color_arr[8] = 8'h0F;
		color_arr[9] = 8'h0F;
		color_arr[10] = 8'h0F;
		color_arr[11] = 8'h0F;
		color_arr[12] = 8'h0F;
		color_arr[13] = 8'h0F;
		color_arr[14] = 8'h0F;
		color_arr[15] = 8'h0F;
		color_arr[16] = 8'h0F;
		color_arr[17] = 8'h0F;
		color_arr[18] = 8'h0F;
		color_arr[19] = 8'h0F;
		color_arr[20] = 8'h0F;
		color_arr[21] = 8'h0F;
		color_arr[22] = 8'h0F;
		color_arr[23] = 8'h0F;
		color_arr[24] = 8'h0F;
		color_arr[25] = 8'h0F;
		color_arr[26] = 8'h0F;
		color_arr[27] = 8'h0F;
		color_arr[28] = 8'h0F;
		color_arr[29] = 8'h0F;
		color_arr[30] = 8'h0F;
		color_arr[31] = 8'h0F;
		color_arr[32] = 8'h0F;
		color_arr[33] = 8'h0F;
		color_arr[34] = 8'h0F;
		color_arr[35] = 8'h0F;
		color_arr[36] = 8'h0F;
		color_arr[37] = 8'h0F;
		color_arr[38] = 8'h0F;
		color_arr[39] = 8'h0F;
		color_arr[40] = 8'h0F;
		color_arr[41] = 8'h0F;
		color_arr[42] = 8'h0F;
		color_arr[43] = 8'h0F;
		color_arr[44] = 8'h0F;
		color_arr[45] = 8'h0F;
		color_arr[46] = 8'h0F;
		color_arr[47] = 8'h0F;
		color_arr[48] = 8'h0F;
		color_arr[49] = 8'h0F;
		color_arr[50] = 8'h0F;
		color_arr[51] = 8'h0F;
		color_arr[52] = 8'h0F;
		color_arr[53] = 8'h0F;
		color_arr[54] = 8'h0F;
		color_arr[55] = 8'h0F;
		color_arr[56] = 8'h0F;
		color_arr[57] = 8'h0F;
		color_arr[58] = 8'h0F;
		color_arr[59] = 8'h0F;
		color_arr[60] = 8'h0F;
		color_arr[61] = 8'h0F;
		color_arr[62] = 8'h0F;
		color_arr[63] = 8'h0F;
		color_arr[64] = 8'h0F;
		color_arr[65] = 8'h0F;
		color_arr[66] = 8'h0F;
		color_arr[67] = 8'h0F;
		color_arr[68] = 8'h0F;
		color_arr[69] = 8'h0F;
		color_arr[70] = 8'h0F;
		color_arr[71] = 8'h0F;
		color_arr[72] = 8'h0F;
		color_arr[73] = 8'h0F;
		color_arr[74] = 8'h0F;
		color_arr[75] = 8'h0F;
		color_arr[76] = 8'h0F;
		color_arr[77] = 8'h0F;
		color_arr[78] = 8'h0F;
		color_arr[79] = 8'h0F;
		color_arr[80] = 8'h0F;
		color_arr[81] = 8'h0F;
		color_arr[82] = 8'h0F;
		color_arr[83] = 8'h0F;
		color_arr[84] = 8'h0F;
		color_arr[85] = 8'h0F;
		color_arr[86] = 8'h0F;
		color_arr[87] = 8'h0F;
		color_arr[88] = 8'h0F;
		color_arr[89] = 8'h0F;
		color_arr[90] = 8'h0F;
		color_arr[91] = 8'h0F;
		color_arr[92] = 8'h0F;
		color_arr[93] = 8'h0F;
		color_arr[94] = 8'h0F;
		color_arr[95] = 8'h0F;
		color_arr[96] = 8'h0F;
		color_arr[97] = 8'h0F;
		color_arr[98] = 8'h0F;
		color_arr[99] = 8'h0F;
		color_arr[100] = 8'h0F;
		color_arr[101] = 8'h0F;
		color_arr[102] = 8'h0F;
		color_arr[103] = 8'h0F;
		color_arr[104] = 8'h0F;
		color_arr[105] = 8'h0F;
		color_arr[106] = 8'h0F;
		color_arr[107] = 8'h0F;
		color_arr[108] = 8'h0F;
		color_arr[109] = 8'h0F;
		color_arr[110] = 8'h0F;
		color_arr[111] = 8'h0F;
		color_arr[112] = 8'h0F;
		color_arr[113] = 8'h0F;
		color_arr[114] = 8'h0F;
		color_arr[115] = 8'h0F;
		color_arr[116] = 8'h0F;
		color_arr[117] = 8'h0F;
		color_arr[118] = 8'h0F;
		color_arr[119] = 8'h0F;
		color_arr[120] = 8'h0F;
		color_arr[121] = 8'h0F;
		color_arr[122] = 8'h0F;
		color_arr[123] = 8'h0F;
		color_arr[124] = 8'h0F;
		color_arr[125] = 8'h0F;
		color_arr[126] = 8'h0F;
		color_arr[127] = 8'h0F;
		color_arr[128] = 8'h0F;
		color_arr[129] = 8'h0F;
		color_arr[130] = 8'h0F;
		color_arr[131] = 8'h0F;
		color_arr[132] = 8'h0F;
		color_arr[133] = 8'h0F;
		color_arr[134] = 8'h0F;
		color_arr[135] = 8'h0F;
		color_arr[136] = 8'h0F;
		color_arr[137] = 8'h0F;
		color_arr[138] = 8'h0F;
		color_arr[139] = 8'h0F;
		color_arr[140] = 8'h0F;
		color_arr[141] = 8'h0F;
		color_arr[142] = 8'h0F;
		color_arr[143] = 8'h0F;
		color_arr[144] = 8'h0F;
		color_arr[145] = 8'h0F;
		color_arr[146] = 8'h0F;
		color_arr[147] = 8'h0F;
		color_arr[148] = 8'h0F;
		color_arr[149] = 8'h0F;
		color_arr[150] = 8'h0F;
		color_arr[151] = 8'h0F;
		color_arr[152] = 8'h0F;
		color_arr[153] = 8'h0F;
		color_arr[154] = 8'h0F;
		color_arr[155] = 8'h0F;
		color_arr[156] = 8'h0F;
		color_arr[157] = 8'h0F;
		color_arr[158] = 8'h0F;
		color_arr[159] = 8'h0F;
		color_arr[160] = 8'h0F;
		color_arr[161] = 8'h0F;
		color_arr[162] = 8'h0F;
		color_arr[163] = 8'h0F;
		color_arr[164] = 8'h0F;
		color_arr[165] = 8'h0F;
		color_arr[166] = 8'h0F;
		color_arr[167] = 8'h0F;
		color_arr[168] = 8'h0F;
		color_arr[169] = 8'h0F;
		color_arr[170] = 8'h0F;
		color_arr[171] = 8'h0F;
		color_arr[172] = 8'h0F;
		color_arr[173] = 8'h0F;
		color_arr[174] = 8'h0F;
		color_arr[175] = 8'h0F;
		color_arr[176] = 8'h0F;
		color_arr[177] = 8'h0F;
		color_arr[178] = 8'h0F;
		color_arr[179] = 8'h0F;
		color_arr[180] = 8'h0F;
		color_arr[181] = 8'h0F;
		color_arr[182] = 8'h0F;
		color_arr[183] = 8'h0F;
		color_arr[184] = 8'h0F;
		color_arr[185] = 8'h0F;
		color_arr[186] = 8'h0F;
		color_arr[187] = 8'h0F;
		color_arr[188] = 8'h0F;
		color_arr[189] = 8'h0F;
		color_arr[190] = 8'h0F;
		color_arr[191] = 8'h0F;
		color_arr[192] = 8'h0F;
		color_arr[193] = 8'h0F;
		color_arr[194] = 8'h0F;
		color_arr[195] = 8'h0F;
		color_arr[196] = 8'h0F;
		color_arr[197] = 8'h0F;
		color_arr[198] = 8'h0F;
		color_arr[199] = 8'h0F;
		color_arr[200] = 8'h0F;
		color_arr[201] = 8'h0F;
		color_arr[202] = 8'h0F;
		color_arr[203] = 8'h0F;
		color_arr[204] = 8'h0F;
		color_arr[205] = 8'h0F;
		color_arr[206] = 8'h0F;
		color_arr[207] = 8'h0F;
		color_arr[208] = 8'h0F;
		color_arr[209] = 8'h0F;
		color_arr[210] = 8'h0F;
		color_arr[211] = 8'h0F;
		color_arr[212] = 8'h0F;
		color_arr[213] = 8'h0F;
		color_arr[214] = 8'h0F;
		color_arr[215] = 8'h0F;
		color_arr[216] = 8'h0F;
		color_arr[217] = 8'h0F;
		color_arr[218] = 8'h0F;
		color_arr[219] = 8'h0F;
		color_arr[220] = 8'h0F;
		color_arr[221] = 8'h0F;
		color_arr[222] = 8'h0F;
		color_arr[223] = 8'h0F;
		color_arr[224] = 8'h0F;
		color_arr[225] = 8'h0F;
		color_arr[226] = 8'h0F;
		color_arr[227] = 8'h0F;
		color_arr[228] = 8'h0F;
		color_arr[229] = 8'h0F;
		color_arr[230] = 8'h0F;
		color_arr[231] = 8'h0F;
		color_arr[232] = 8'h0F;
		color_arr[233] = 8'h0F;
		color_arr[234] = 8'h0F;
		color_arr[235] = 8'h0F;
		color_arr[236] = 8'h0F;
		color_arr[237] = 8'h0F;
		color_arr[238] = 8'h0F;
		color_arr[239] = 8'h0F;
		color_arr[240] = 8'h0F;
		color_arr[241] = 8'h0F;
		color_arr[242] = 8'h0F;
		color_arr[243] = 8'h0F;
		color_arr[244] = 8'h0F;
		color_arr[245] = 8'h0F;
		color_arr[246] = 8'h0F;
		color_arr[247] = 8'h0F;
		color_arr[248] = 8'h0F;
		color_arr[249] = 8'h0F;
		color_arr[250] = 8'h0F;
		color_arr[251] = 8'h0F;
		color_arr[252] = 8'h0F;
		color_arr[253] = 8'h0F;
		color_arr[254] = 8'h0F;
		color_arr[255] = 8'h0F;
		color_arr[256] = 8'h0F;
		color_arr[257] = 8'h0F;
		color_arr[258] = 8'h0F;
		color_arr[259] = 8'h0F;
		color_arr[260] = 8'h0F;
		color_arr[261] = 8'h0F;
		color_arr[262] = 8'h0F;
		color_arr[263] = 8'h0F;
		color_arr[264] = 8'h0F;
		color_arr[265] = 8'h0F;
		color_arr[266] = 8'h0F;
		color_arr[267] = 8'h0F;
		color_arr[268] = 8'h0F;
		color_arr[269] = 8'h0F;
		color_arr[270] = 8'h0F;
		color_arr[271] = 8'h0F;
		color_arr[272] = 8'h0F;
		color_arr[273] = 8'h0F;
		color_arr[274] = 8'h0F;
		color_arr[275] = 8'h0F;
		color_arr[276] = 8'h0F;
		color_arr[277] = 8'h0F;
		color_arr[278] = 8'h0F;
		color_arr[279] = 8'h0F;
		color_arr[280] = 8'h0F;
		color_arr[281] = 8'h0F;
		color_arr[282] = 8'h0F;
		color_arr[283] = 8'h0F;
		color_arr[284] = 8'h0F;
		color_arr[285] = 8'h0F;
		color_arr[286] = 8'h0F;
		color_arr[287] = 8'h0F;
		color_arr[288] = 8'h0F;
		color_arr[289] = 8'h0F;
		color_arr[290] = 8'h0F;
		color_arr[291] = 8'h0F;
		color_arr[292] = 8'h0F;
		color_arr[293] = 8'h0F;
		color_arr[294] = 8'h0F;
		color_arr[295] = 8'h0F;
		color_arr[296] = 8'h0F;
		color_arr[297] = 8'h0F;
		color_arr[298] = 8'h0F;
		color_arr[299] = 8'h0F;
		color_arr[300] = 8'h0F;
		color_arr[301] = 8'h0F;
		color_arr[302] = 8'h0F;
		color_arr[303] = 8'h0F;
		color_arr[304] = 8'h0F;
		color_arr[305] = 8'h0F;
		color_arr[306] = 8'h0F;
		color_arr[307] = 8'h0F;
		color_arr[308] = 8'h0F;
		color_arr[309] = 8'h0F;
		color_arr[310] = 8'h0F;
		color_arr[311] = 8'h0F;
		color_arr[312] = 8'h0F;
		color_arr[313] = 8'h0F;
		color_arr[314] = 8'h0F;
		color_arr[315] = 8'h0F;
		color_arr[316] = 8'h0F;
		color_arr[317] = 8'h0F;
		color_arr[318] = 8'h0F;
		color_arr[319] = 8'h0F;
		color_arr[320] = 8'h0F;
		color_arr[321] = 8'h0F;
		color_arr[322] = 8'h0F;
		color_arr[323] = 8'h0F;
		color_arr[324] = 8'h0F;
		color_arr[325] = 8'h0F;
		color_arr[326] = 8'h0F;
		color_arr[327] = 8'h0F;
		color_arr[328] = 8'h0F;
		color_arr[329] = 8'h0F;
		color_arr[330] = 8'h0F;
		color_arr[331] = 8'h0F;
		color_arr[332] = 8'h0F;
		color_arr[333] = 8'h0F;
		color_arr[334] = 8'h0F;
		color_arr[335] = 8'h0F;
		color_arr[336] = 8'h0F;
		color_arr[337] = 8'h0F;
		color_arr[338] = 8'h0F;
		color_arr[339] = 8'h0F;
		color_arr[340] = 8'h0F;
		color_arr[341] = 8'h0F;
		color_arr[342] = 8'h0F;
		color_arr[343] = 8'h0F;
		color_arr[344] = 8'h0F;
		color_arr[345] = 8'h0F;
		color_arr[346] = 8'h0F;
		color_arr[347] = 8'h0F;
		color_arr[348] = 8'h0F;
		color_arr[349] = 8'h0F;
		color_arr[350] = 8'h0F;
		color_arr[351] = 8'h0F;
		color_arr[352] = 8'h0F;
		color_arr[353] = 8'h0F;
		color_arr[354] = 8'h0F;
		color_arr[355] = 8'h0F;
		color_arr[356] = 8'h0F;
		color_arr[357] = 8'h0F;
		color_arr[358] = 8'h0F;
		color_arr[359] = 8'h0F;
		color_arr[360] = 8'h0F;
		color_arr[361] = 8'h0F;
		color_arr[362] = 8'h0F;
		color_arr[363] = 8'h0F;
		color_arr[364] = 8'h0F;
		color_arr[365] = 8'h0F;
		color_arr[366] = 8'h0F;
		color_arr[367] = 8'h0F;
		color_arr[368] = 8'h0F;
		color_arr[369] = 8'h0F;
		color_arr[370] = 8'h0F;
		color_arr[371] = 8'h0F;
		color_arr[372] = 8'h0F;
		color_arr[373] = 8'h0F;
		color_arr[374] = 8'h0F;
		color_arr[375] = 8'h0F;
		color_arr[376] = 8'h0F;
		color_arr[377] = 8'h0F;
		color_arr[378] = 8'h0F;
		color_arr[379] = 8'h0F;
		color_arr[380] = 8'h0F;
		color_arr[381] = 8'h0F;
		color_arr[382] = 8'h0F;
		color_arr[383] = 8'h0F;
		color_arr[384] = 8'h0F;
		color_arr[385] = 8'h0F;
		color_arr[386] = 8'h0F;
		color_arr[387] = 8'h0F;
		color_arr[388] = 8'h0F;
		color_arr[389] = 8'h0F;
		color_arr[390] = 8'h0F;
		color_arr[391] = 8'h0F;
		color_arr[392] = 8'h0F;
		color_arr[393] = 8'h0F;
		color_arr[394] = 8'h0F;
		color_arr[395] = 8'h0F;
		color_arr[396] = 8'h0F;
		color_arr[397] = 8'h0F;
		color_arr[398] = 8'h0F;
		color_arr[399] = 8'h0F;
		color_arr[400] = 8'h0F;
		color_arr[401] = 8'h0F;
		color_arr[402] = 8'h0F;
		color_arr[403] = 8'h0F;
		color_arr[404] = 8'h0F;
		color_arr[405] = 8'h0F;
		color_arr[406] = 8'h0F;
		color_arr[407] = 8'h0F;
		color_arr[408] = 8'h0F;
		color_arr[409] = 8'h0F;
		color_arr[410] = 8'h0F;
		color_arr[411] = 8'h0F;
		color_arr[412] = 8'h0F;
		color_arr[413] = 8'h0F;
		color_arr[414] = 8'h0F;
		color_arr[415] = 8'h0F;
		color_arr[416] = 8'h0F;
		color_arr[417] = 8'h0F;
		color_arr[418] = 8'h0F;
		color_arr[419] = 8'h0F;
		color_arr[420] = 8'h0F;
		color_arr[421] = 8'h0F;
		color_arr[422] = 8'h0F;
		color_arr[423] = 8'h0F;
		color_arr[424] = 8'h0F;
		color_arr[425] = 8'h0F;
		color_arr[426] = 8'h0F;
		color_arr[427] = 8'h0F;
		color_arr[428] = 8'h0F;
		color_arr[429] = 8'h0F;
		color_arr[430] = 8'h0F;
		color_arr[431] = 8'h0F;
		color_arr[432] = 8'h0F;
		color_arr[433] = 8'h0F;
		color_arr[434] = 8'h0F;
		color_arr[435] = 8'h0F;
		color_arr[436] = 8'h0F;
		color_arr[437] = 8'h0F;
		color_arr[438] = 8'h0F;
		color_arr[439] = 8'h0F;
		color_arr[440] = 8'h0F;
		color_arr[441] = 8'h0F;
		color_arr[442] = 8'h0F;
		color_arr[443] = 8'h0F;
		color_arr[444] = 8'h0F;
		color_arr[445] = 8'h0F;
		color_arr[446] = 8'h0F;
		color_arr[447] = 8'h0F;
		color_arr[448] = 8'h0F;
		color_arr[449] = 8'h0F;
		color_arr[450] = 8'h0F;
		color_arr[451] = 8'h0F;
		color_arr[452] = 8'h0F;
		color_arr[453] = 8'h0F;
		color_arr[454] = 8'h0F;
		color_arr[455] = 8'h0F;
		color_arr[456] = 8'h0F;
		color_arr[457] = 8'h0F;
		color_arr[458] = 8'h0F;
		color_arr[459] = 8'h0F;
		color_arr[460] = 8'h0F;
		color_arr[461] = 8'h0F;
		color_arr[462] = 8'h0F;
		color_arr[463] = 8'h0F;
		color_arr[464] = 8'h0F;
		color_arr[465] = 8'h0F;
		color_arr[466] = 8'h0F;
		color_arr[467] = 8'h0F;
		color_arr[468] = 8'h0F;
		color_arr[469] = 8'h0F;
		color_arr[470] = 8'h0F;
		color_arr[471] = 8'h0F;
		color_arr[472] = 8'h0F;
		color_arr[473] = 8'h0F;
		color_arr[474] = 8'h0F;
		color_arr[475] = 8'h0F;
		color_arr[476] = 8'h0F;
		color_arr[477] = 8'h0F;
		color_arr[478] = 8'h0F;
		color_arr[479] = 8'h0F;
		color_arr[480] = 8'h0F;
		color_arr[481] = 8'h0F;
		color_arr[482] = 8'h0F;
		color_arr[483] = 8'h0F;
		color_arr[484] = 8'h0F;
		color_arr[485] = 8'h0F;
		color_arr[486] = 8'h0F;
		color_arr[487] = 8'h0F;
		color_arr[488] = 8'h0F;
		color_arr[489] = 8'h0F;
		color_arr[490] = 8'h0F;
		color_arr[491] = 8'h0F;
		color_arr[492] = 8'h0F;
		color_arr[493] = 8'h0F;
		color_arr[494] = 8'h0F;
		color_arr[495] = 8'h0F;
		color_arr[496] = 8'h0F;
		color_arr[497] = 8'h0F;
		color_arr[498] = 8'h0F;
		color_arr[499] = 8'h0F;
		color_arr[500] = 8'h0F;
		color_arr[501] = 8'h0F;
		color_arr[502] = 8'h0F;
		color_arr[503] = 8'h0F;
		color_arr[504] = 8'h0F;
		color_arr[505] = 8'h0F;
		color_arr[506] = 8'h0F;
		color_arr[507] = 8'h0F;
		color_arr[508] = 8'h0F;
		color_arr[509] = 8'h0F;
		color_arr[510] = 8'h0F;
		color_arr[511] = 8'h0F;
		color_arr[512] = 8'h0F;
		color_arr[513] = 8'h0F;
		color_arr[514] = 8'h0F;
		color_arr[515] = 8'h0F;
		color_arr[516] = 8'h0F;
		color_arr[517] = 8'h0F;
		color_arr[518] = 8'h0F;
		color_arr[519] = 8'h0F;
		color_arr[520] = 8'h0F;
		color_arr[521] = 8'h0F;
		color_arr[522] = 8'h0F;
		color_arr[523] = 8'h0F;
		color_arr[524] = 8'h0F;
		color_arr[525] = 8'h0F;
		color_arr[526] = 8'h0F;
		color_arr[527] = 8'h0F;
		color_arr[528] = 8'h0F;
		color_arr[529] = 8'h0F;
		color_arr[530] = 8'h0F;
		color_arr[531] = 8'h0F;
		color_arr[532] = 8'h0F;
		color_arr[533] = 8'h0F;
		color_arr[534] = 8'h0F;
		color_arr[535] = 8'h0F;
		color_arr[536] = 8'h0F;
		color_arr[537] = 8'h0F;
		color_arr[538] = 8'h0F;
		color_arr[539] = 8'h0F;
		color_arr[540] = 8'h0F;
		color_arr[541] = 8'h0F;
		color_arr[542] = 8'h0F;
		color_arr[543] = 8'h0F;
		color_arr[544] = 8'h0F;
		color_arr[545] = 8'h0F;
		color_arr[546] = 8'h0F;
		color_arr[547] = 8'h0F;
		color_arr[548] = 8'h0F;
		color_arr[549] = 8'h0F;
		color_arr[550] = 8'h0F;
		color_arr[551] = 8'h0F;
		color_arr[552] = 8'h0F;
		color_arr[553] = 8'h0F;
		color_arr[554] = 8'h0F;
		color_arr[555] = 8'h0F;
		color_arr[556] = 8'h0F;
		color_arr[557] = 8'h0F;
		color_arr[558] = 8'h0F;
		color_arr[559] = 8'h0F;
		color_arr[560] = 8'h0F;
		color_arr[561] = 8'h0F;
		color_arr[562] = 8'h0F;
		color_arr[563] = 8'h0F;
		color_arr[564] = 8'h0F;
		color_arr[565] = 8'h0F;
		color_arr[566] = 8'h0F;
		color_arr[567] = 8'h0F;
		color_arr[568] = 8'h0F;
		color_arr[569] = 8'h0F;
		color_arr[570] = 8'h0F;
		color_arr[571] = 8'h0F;
		color_arr[572] = 8'h0F;
		color_arr[573] = 8'h0F;
		color_arr[574] = 8'h0F;
		color_arr[575] = 8'h0F;
		color_arr[576] = 8'h0F;
		color_arr[577] = 8'h0F;
		color_arr[578] = 8'h0F;
		color_arr[579] = 8'h0F;
		color_arr[580] = 8'h0F;
		color_arr[581] = 8'h0F;
		color_arr[582] = 8'h0F;
		color_arr[583] = 8'h0F;
		color_arr[584] = 8'h0F;
		color_arr[585] = 8'h0F;
		color_arr[586] = 8'h0F;
		color_arr[587] = 8'h0F;
		color_arr[588] = 8'h0F;
		color_arr[589] = 8'h0F;
		color_arr[590] = 8'h0F;
		color_arr[591] = 8'h0F;
		color_arr[592] = 8'h0F;
		color_arr[593] = 8'h0F;
		color_arr[594] = 8'h0F;
		color_arr[595] = 8'h0F;
		color_arr[596] = 8'h0F;
		color_arr[597] = 8'h0F;
		color_arr[598] = 8'h0F;
		color_arr[599] = 8'h0F;
		color_arr[600] = 8'h0F;
		color_arr[601] = 8'h0F;
		color_arr[602] = 8'h0F;
		color_arr[603] = 8'h0F;
		color_arr[604] = 8'h0F;
		color_arr[605] = 8'h0F;
		color_arr[606] = 8'h0F;
		color_arr[607] = 8'h0F;
		color_arr[608] = 8'h0F;
		color_arr[609] = 8'h0F;
		color_arr[610] = 8'h0F;
		color_arr[611] = 8'h0F;
		color_arr[612] = 8'h0F;
		color_arr[613] = 8'h0F;
		color_arr[614] = 8'h0F;
		color_arr[615] = 8'h0F;
		color_arr[616] = 8'h0F;
		color_arr[617] = 8'h0F;
		color_arr[618] = 8'h0F;
		color_arr[619] = 8'h0F;
		color_arr[620] = 8'h0F;
		color_arr[621] = 8'h0F;
		color_arr[622] = 8'h0F;
		color_arr[623] = 8'h0F;
		color_arr[624] = 8'h0F;
		color_arr[625] = 8'h0F;
		color_arr[626] = 8'h0F;
		color_arr[627] = 8'h0F;
		color_arr[628] = 8'h0F;
		color_arr[629] = 8'h0F;
		color_arr[630] = 8'h0F;
		color_arr[631] = 8'h0F;
		color_arr[632] = 8'h0F;
		color_arr[633] = 8'h0F;
		color_arr[634] = 8'h0F;
		color_arr[635] = 8'h0F;
		color_arr[636] = 8'h0F;
		color_arr[637] = 8'h0F;
		color_arr[638] = 8'h0F;
		color_arr[639] = 8'h0F;
		color_arr[640] = 8'h0F;
		color_arr[641] = 8'h0F;
		color_arr[642] = 8'h0F;
		color_arr[643] = 8'h0F;
		color_arr[644] = 8'h0F;
		color_arr[645] = 8'h0F;
		color_arr[646] = 8'h0F;
		color_arr[647] = 8'h0F;
		color_arr[648] = 8'h0F;
		color_arr[649] = 8'h0F;
		color_arr[650] = 8'h0F;
		color_arr[651] = 8'h0F;
		color_arr[652] = 8'h0F;
		color_arr[653] = 8'h0F;
		color_arr[654] = 8'h0F;
		color_arr[655] = 8'h0F;
		color_arr[656] = 8'h0F;
		color_arr[657] = 8'h0F;
		color_arr[658] = 8'h0F;
		color_arr[659] = 8'h0F;
		color_arr[660] = 8'h0F;
		color_arr[661] = 8'h0F;
		color_arr[662] = 8'h0F;
		color_arr[663] = 8'h0F;
		color_arr[664] = 8'h0F;
		color_arr[665] = 8'h0F;
		color_arr[666] = 8'h0F;
		color_arr[667] = 8'h0F;
		color_arr[668] = 8'h0F;
		color_arr[669] = 8'h0F;
		color_arr[670] = 8'h0F;
		color_arr[671] = 8'h0F;
		color_arr[672] = 8'h0F;
		color_arr[673] = 8'h0F;
		color_arr[674] = 8'h0F;
		color_arr[675] = 8'h0F;
		color_arr[676] = 8'h0F;
		color_arr[677] = 8'h0F;
		color_arr[678] = 8'h0F;
		color_arr[679] = 8'h0F;
		color_arr[680] = 8'h0F;
		color_arr[681] = 8'h0F;
		color_arr[682] = 8'h0F;
		color_arr[683] = 8'h0F;
		color_arr[684] = 8'h0F;
		color_arr[685] = 8'h0F;
		color_arr[686] = 8'h0F;
		color_arr[687] = 8'h0F;
		color_arr[688] = 8'h0F;
		color_arr[689] = 8'h0F;
		color_arr[690] = 8'h0F;
		color_arr[691] = 8'h0F;
		color_arr[692] = 8'h0F;
		color_arr[693] = 8'h0F;
		color_arr[694] = 8'h0F;
		color_arr[695] = 8'h0F;
		color_arr[696] = 8'h0F;
		color_arr[697] = 8'h0F;
		color_arr[698] = 8'h0F;
		color_arr[699] = 8'h0F;
		color_arr[700] = 8'h0F;
		color_arr[701] = 8'h0F;
		color_arr[702] = 8'h0F;
		color_arr[703] = 8'h0F;
		color_arr[704] = 8'h0F;
		color_arr[705] = 8'h0F;
		color_arr[706] = 8'h0F;
		color_arr[707] = 8'h0F;
		color_arr[708] = 8'h0F;
		color_arr[709] = 8'h0F;
		color_arr[710] = 8'h0F;
		color_arr[711] = 8'h0F;
		color_arr[712] = 8'h0F;
		color_arr[713] = 8'h0F;
		color_arr[714] = 8'h0F;
		color_arr[715] = 8'h0F;
		color_arr[716] = 8'h0F;
		color_arr[717] = 8'h0F;
		color_arr[718] = 8'h0F;
		color_arr[719] = 8'h0F;
		color_arr[720] = 8'h0F;
		color_arr[721] = 8'h0F;
		color_arr[722] = 8'h0F;
		color_arr[723] = 8'h0F;
		color_arr[724] = 8'h0F;
		color_arr[725] = 8'h0F;
		color_arr[726] = 8'h0F;
		color_arr[727] = 8'h0F;
		color_arr[728] = 8'h0F;
		color_arr[729] = 8'h0F;
		color_arr[730] = 8'h0F;
		color_arr[731] = 8'h0F;
		color_arr[732] = 8'h0F;
		color_arr[733] = 8'h0F;
		color_arr[734] = 8'h0F;
		color_arr[735] = 8'h0F;
		color_arr[736] = 8'h0F;
		color_arr[737] = 8'h0F;
		color_arr[738] = 8'h0F;
		color_arr[739] = 8'h0F;
		color_arr[740] = 8'h0F;
		color_arr[741] = 8'h0F;
		color_arr[742] = 8'h0F;
		color_arr[743] = 8'h0F;
		color_arr[744] = 8'h0F;
		color_arr[745] = 8'h0F;
		color_arr[746] = 8'h0F;
		color_arr[747] = 8'h0F;
		color_arr[748] = 8'h0F;
		color_arr[749] = 8'h0F;
		color_arr[750] = 8'h0F;
		color_arr[751] = 8'h0F;
		color_arr[752] = 8'h0F;
		color_arr[753] = 8'h0F;
		color_arr[754] = 8'h0F;
		color_arr[755] = 8'h0F;
		color_arr[756] = 8'h0F;
		color_arr[757] = 8'h0F;
		color_arr[758] = 8'h0F;
		color_arr[759] = 8'h0F;
		color_arr[760] = 8'h0F;
		color_arr[761] = 8'h0F;
		color_arr[762] = 8'h0F;
		color_arr[763] = 8'h0F;
		color_arr[764] = 8'h0F;
		color_arr[765] = 8'h0F;
		color_arr[766] = 8'h0F;
		color_arr[767] = 8'h0F;
		color_arr[768] = 8'h0F;
		color_arr[769] = 8'h0F;
		color_arr[770] = 8'h0F;
		color_arr[771] = 8'h0F;
		color_arr[772] = 8'h0F;
		color_arr[773] = 8'h0F;
		color_arr[774] = 8'h0F;
		color_arr[775] = 8'h0F;
		color_arr[776] = 8'h0F;
		color_arr[777] = 8'h0F;
		color_arr[778] = 8'h0F;
		color_arr[779] = 8'h0F;
		color_arr[780] = 8'h0F;
		color_arr[781] = 8'h0F;
		color_arr[782] = 8'h0F;
		color_arr[783] = 8'h0F;
		color_arr[784] = 8'h0F;
		color_arr[785] = 8'h0F;
		color_arr[786] = 8'h0F;
		color_arr[787] = 8'h0F;
		color_arr[788] = 8'h0F;
		color_arr[789] = 8'h0F;
		color_arr[790] = 8'h0F;
		color_arr[791] = 8'h0F;
		color_arr[792] = 8'h0F;
		color_arr[793] = 8'h0F;
		color_arr[794] = 8'h0F;
		color_arr[795] = 8'h0F;
		color_arr[796] = 8'h0F;
		color_arr[797] = 8'h0F;
		color_arr[798] = 8'h0F;
		color_arr[799] = 8'h0F;
		color_arr[800] = 8'h0F;
		color_arr[801] = 8'h0F;
		color_arr[802] = 8'h0F;
		color_arr[803] = 8'h0F;
		color_arr[804] = 8'h0F;
		color_arr[805] = 8'h0F;
		color_arr[806] = 8'h0F;
		color_arr[807] = 8'h0F;
		color_arr[808] = 8'h0F;
		color_arr[809] = 8'h0F;
		color_arr[810] = 8'h0F;
		color_arr[811] = 8'h0F;
		color_arr[812] = 8'h0F;
		color_arr[813] = 8'h0F;
		color_arr[814] = 8'h0F;
		color_arr[815] = 8'h0F;
		color_arr[816] = 8'h0F;
		color_arr[817] = 8'h0F;
		color_arr[818] = 8'h0F;
		color_arr[819] = 8'h0F;
		color_arr[820] = 8'h0F;
		color_arr[821] = 8'h0F;
		color_arr[822] = 8'h0F;
		color_arr[823] = 8'h0F;
		color_arr[824] = 8'h0F;
		color_arr[825] = 8'h0F;
		color_arr[826] = 8'h0F;
		color_arr[827] = 8'h0F;
		color_arr[828] = 8'h0F;
		color_arr[829] = 8'h0F;
		color_arr[830] = 8'h0F;
		color_arr[831] = 8'h0F;
		color_arr[832] = 8'h0F;
		color_arr[833] = 8'h0F;
		color_arr[834] = 8'h0F;
		color_arr[835] = 8'h0F;
		color_arr[836] = 8'h0F;
		color_arr[837] = 8'h0F;
		color_arr[838] = 8'h0F;
		color_arr[839] = 8'h0F;
		color_arr[840] = 8'h0F;
		color_arr[841] = 8'h0F;
		color_arr[842] = 8'h0F;
		color_arr[843] = 8'h0F;
		color_arr[844] = 8'h0F;
		color_arr[845] = 8'h0F;
		color_arr[846] = 8'h0F;
		color_arr[847] = 8'h0F;
		color_arr[848] = 8'h0F;
		color_arr[849] = 8'h0F;
		color_arr[850] = 8'h0F;
		color_arr[851] = 8'h0F;
		color_arr[852] = 8'h0F;
		color_arr[853] = 8'h0F;
		color_arr[854] = 8'h0F;
		color_arr[855] = 8'h0F;
		color_arr[856] = 8'h0F;
		color_arr[857] = 8'h0F;
		color_arr[858] = 8'h0F;
		color_arr[859] = 8'h0F;
		color_arr[860] = 8'h0F;
		color_arr[861] = 8'h0F;
		color_arr[862] = 8'h0F;
		color_arr[863] = 8'h0F;
		color_arr[864] = 8'h0F;
		color_arr[865] = 8'h0F;
		color_arr[866] = 8'h0F;
		color_arr[867] = 8'h0F;
		color_arr[868] = 8'h0F;
		color_arr[869] = 8'h0F;
		color_arr[870] = 8'h0F;
		color_arr[871] = 8'h0F;
		color_arr[872] = 8'h0F;
		color_arr[873] = 8'h0F;
		color_arr[874] = 8'h0F;
		color_arr[875] = 8'h0F;
		color_arr[876] = 8'h0F;
		color_arr[877] = 8'h0F;
		color_arr[878] = 8'h0F;
		color_arr[879] = 8'h0F;
		color_arr[880] = 8'h0F;
		color_arr[881] = 8'h0F;
		color_arr[882] = 8'h0F;
		color_arr[883] = 8'h0F;
		color_arr[884] = 8'h0F;
		color_arr[885] = 8'h0F;
		color_arr[886] = 8'h0F;
		color_arr[887] = 8'h0F;
		color_arr[888] = 8'h0F;
		color_arr[889] = 8'h0F;
		color_arr[890] = 8'h0F;
		color_arr[891] = 8'h0F;
		color_arr[892] = 8'h0F;
		color_arr[893] = 8'h0F;
		color_arr[894] = 8'h0F;
		color_arr[895] = 8'h0F;
		color_arr[896] = 8'h0F;
		color_arr[897] = 8'h0F;
		color_arr[898] = 8'h0F;
		color_arr[899] = 8'h0F;
		color_arr[900] = 8'h0F;
		color_arr[901] = 8'h0F;
		color_arr[902] = 8'h0F;
		color_arr[903] = 8'h0F;
		color_arr[904] = 8'h0F;
		color_arr[905] = 8'h0F;
		color_arr[906] = 8'h0F;
		color_arr[907] = 8'h0F;
		color_arr[908] = 8'h0F;
		color_arr[909] = 8'h0F;
		color_arr[910] = 8'h0F;
		color_arr[911] = 8'h0F;
		color_arr[912] = 8'h0F;
		color_arr[913] = 8'h0F;
		color_arr[914] = 8'h0F;
		color_arr[915] = 8'h0F;
		color_arr[916] = 8'h0F;
		color_arr[917] = 8'h0F;
		color_arr[918] = 8'h0F;
		color_arr[919] = 8'h0F;
		color_arr[920] = 8'h0F;
		color_arr[921] = 8'h0F;
		color_arr[922] = 8'h0F;
		color_arr[923] = 8'h0F;
		color_arr[924] = 8'h0F;
		color_arr[925] = 8'h0F;
		color_arr[926] = 8'h0F;
		color_arr[927] = 8'h0F;
		color_arr[928] = 8'h0F;
		color_arr[929] = 8'h0F;
		color_arr[930] = 8'h0F;
		color_arr[931] = 8'h0F;
		color_arr[932] = 8'h0F;
		color_arr[933] = 8'h0F;
		color_arr[934] = 8'h0F;
		color_arr[935] = 8'h0F;
		color_arr[936] = 8'h0F;
		color_arr[937] = 8'h0F;
		color_arr[938] = 8'h0F;
		color_arr[939] = 8'h0F;
		color_arr[940] = 8'h0F;
		color_arr[941] = 8'h0F;
		color_arr[942] = 8'h0F;
		color_arr[943] = 8'h0F;
		color_arr[944] = 8'h0F;
		color_arr[945] = 8'h0F;
		color_arr[946] = 8'h0F;
		color_arr[947] = 8'h0F;
		color_arr[948] = 8'h0F;
		color_arr[949] = 8'h0F;
		color_arr[950] = 8'h0F;
		color_arr[951] = 8'h0F;
		color_arr[952] = 8'h0F;
		color_arr[953] = 8'h0F;
		color_arr[954] = 8'h0F;
		color_arr[955] = 8'h0F;
		color_arr[956] = 8'h0F;
		color_arr[957] = 8'h0F;
		color_arr[958] = 8'h0F;
		color_arr[959] = 8'h0F;
		color_arr[960] = 8'h0F;
		color_arr[961] = 8'h0F;
		color_arr[962] = 8'h0F;
		color_arr[963] = 8'h0F;
		color_arr[964] = 8'h0F;
		color_arr[965] = 8'h0F;
		color_arr[966] = 8'h0F;
		color_arr[967] = 8'h0F;
		color_arr[968] = 8'h0F;
		color_arr[969] = 8'h0F;
		color_arr[970] = 8'h0F;
		color_arr[971] = 8'h0F;
		color_arr[972] = 8'h0F;
		color_arr[973] = 8'h0F;
		color_arr[974] = 8'h0F;
		color_arr[975] = 8'h0F;
		color_arr[976] = 8'h0F;
		color_arr[977] = 8'h0F;
		color_arr[978] = 8'h0F;
		color_arr[979] = 8'h0F;
		color_arr[980] = 8'h0F;
		color_arr[981] = 8'h0F;
		color_arr[982] = 8'h0F;
		color_arr[983] = 8'h0F;
		color_arr[984] = 8'h0F;
		color_arr[985] = 8'h0F;
		color_arr[986] = 8'h0F;
		color_arr[987] = 8'h0F;
		color_arr[988] = 8'h0F;
		color_arr[989] = 8'h0F;
		color_arr[990] = 8'h0F;
		color_arr[991] = 8'h0F;
		color_arr[992] = 8'h0F;
		color_arr[993] = 8'h0F;
		color_arr[994] = 8'h0F;
		color_arr[995] = 8'h0F;
		color_arr[996] = 8'h0F;
		color_arr[997] = 8'h0F;
		color_arr[998] = 8'h0F;
		color_arr[999] = 8'h0F;
		color_arr[1000] = 8'h0F;
		color_arr[1001] = 8'h0F;
		color_arr[1002] = 8'h0F;
		color_arr[1003] = 8'h0F;
		color_arr[1004] = 8'h0F;
		color_arr[1005] = 8'h0F;
		color_arr[1006] = 8'h0F;
		color_arr[1007] = 8'h0F;
		color_arr[1008] = 8'h0F;
		color_arr[1009] = 8'h0F;
		color_arr[1010] = 8'h0F;
		color_arr[1011] = 8'h0F;
		color_arr[1012] = 8'h0F;
		color_arr[1013] = 8'h0F;
		color_arr[1014] = 8'h0F;
		color_arr[1015] = 8'h0F;
		color_arr[1016] = 8'h0F;
		color_arr[1017] = 8'h0F;
		color_arr[1018] = 8'h0F;
		color_arr[1019] = 8'h0F;
		color_arr[1020] = 8'h0F;
		color_arr[1021] = 8'h0F;
		color_arr[1022] = 8'h0F;
		color_arr[1023] = 8'h0F;
		color_arr[1024] = 8'h0F;
		color_arr[1025] = 8'h0F;
		color_arr[1026] = 8'h0F;
		color_arr[1027] = 8'h0F;
		color_arr[1028] = 8'h0F;
		color_arr[1029] = 8'h0F;
		color_arr[1030] = 8'h0F;
		color_arr[1031] = 8'h0F;
		color_arr[1032] = 8'h0F;
		color_arr[1033] = 8'h0F;
		color_arr[1034] = 8'h0F;
		color_arr[1035] = 8'h0F;
		color_arr[1036] = 8'h0F;
		color_arr[1037] = 8'h0F;
		color_arr[1038] = 8'h0F;
		color_arr[1039] = 8'h0F;
		color_arr[1040] = 8'h0F;
		color_arr[1041] = 8'h0F;
		color_arr[1042] = 8'h0F;
		color_arr[1043] = 8'h0F;
		color_arr[1044] = 8'h0F;
		color_arr[1045] = 8'h0F;
		color_arr[1046] = 8'h0F;
		color_arr[1047] = 8'h0F;
		color_arr[1048] = 8'h0F;
		color_arr[1049] = 8'h0F;
		color_arr[1050] = 8'h0F;
		color_arr[1051] = 8'h0F;
		color_arr[1052] = 8'h0F;
		color_arr[1053] = 8'h0F;
		color_arr[1054] = 8'h0F;
		color_arr[1055] = 8'h0F;
		color_arr[1056] = 8'h0F;
		color_arr[1057] = 8'h0F;
		color_arr[1058] = 8'h0F;
		color_arr[1059] = 8'h0F;
		color_arr[1060] = 8'h0F;
		color_arr[1061] = 8'h0F;
		color_arr[1062] = 8'h0F;
		color_arr[1063] = 8'h0F;
		color_arr[1064] = 8'h0F;
		color_arr[1065] = 8'h0F;
		color_arr[1066] = 8'h0F;
		color_arr[1067] = 8'h0F;
		color_arr[1068] = 8'h0F;
		color_arr[1069] = 8'h0F;
		color_arr[1070] = 8'h0F;
		color_arr[1071] = 8'h0F;
		color_arr[1072] = 8'h0F;
		color_arr[1073] = 8'h0F;
		color_arr[1074] = 8'h0F;
		color_arr[1075] = 8'h0F;
		color_arr[1076] = 8'h0F;
		color_arr[1077] = 8'h0F;
		color_arr[1078] = 8'h0F;
		color_arr[1079] = 8'h0F;
		color_arr[1080] = 8'h0F;
		color_arr[1081] = 8'h0F;
		color_arr[1082] = 8'h0F;
		color_arr[1083] = 8'h0F;
		color_arr[1084] = 8'h0F;
		color_arr[1085] = 8'h0F;
		color_arr[1086] = 8'h0F;
		color_arr[1087] = 8'h0F;
		color_arr[1088] = 8'h0F;
		color_arr[1089] = 8'h0F;
		color_arr[1090] = 8'h0F;
		color_arr[1091] = 8'h0F;
		color_arr[1092] = 8'h0F;
		color_arr[1093] = 8'h0F;
		color_arr[1094] = 8'h0F;
		color_arr[1095] = 8'h0F;
		color_arr[1096] = 8'h0F;
		color_arr[1097] = 8'h0F;
		color_arr[1098] = 8'h0F;
		color_arr[1099] = 8'h0F;
		color_arr[1100] = 8'h0F;
		color_arr[1101] = 8'h0F;
		color_arr[1102] = 8'h0F;
		color_arr[1103] = 8'h0F;
		color_arr[1104] = 8'h0F;
		color_arr[1105] = 8'h0F;
		color_arr[1106] = 8'h0F;
		color_arr[1107] = 8'h0F;
		color_arr[1108] = 8'h0F;
		color_arr[1109] = 8'h0F;
		color_arr[1110] = 8'h0F;
		color_arr[1111] = 8'h0F;
		color_arr[1112] = 8'h0F;
		color_arr[1113] = 8'h0F;
		color_arr[1114] = 8'h0F;
		color_arr[1115] = 8'h0F;
		color_arr[1116] = 8'h0F;
		color_arr[1117] = 8'h0F;
		color_arr[1118] = 8'h0F;
		color_arr[1119] = 8'h0F;
		color_arr[1120] = 8'h0F;
		color_arr[1121] = 8'h0F;
		color_arr[1122] = 8'h0F;
		color_arr[1123] = 8'h0F;
		color_arr[1124] = 8'h0F;
		color_arr[1125] = 8'h0F;
		color_arr[1126] = 8'h0F;
		color_arr[1127] = 8'h0F;
		color_arr[1128] = 8'h0F;
		color_arr[1129] = 8'h0F;
		color_arr[1130] = 8'h0F;
		color_arr[1131] = 8'h0F;
		color_arr[1132] = 8'h0F;
		color_arr[1133] = 8'h0F;
		color_arr[1134] = 8'h0F;
		color_arr[1135] = 8'h0F;
		color_arr[1136] = 8'h0F;
		color_arr[1137] = 8'h0F;
		color_arr[1138] = 8'h0F;
		color_arr[1139] = 8'h0F;
		color_arr[1140] = 8'h0F;
		color_arr[1141] = 8'h0F;
		color_arr[1142] = 8'h0F;
		color_arr[1143] = 8'h0F;
		color_arr[1144] = 8'h0F;
		color_arr[1145] = 8'h0F;
		color_arr[1146] = 8'h0F;
		color_arr[1147] = 8'h0F;
		color_arr[1148] = 8'h0F;
		color_arr[1149] = 8'h0F;
		color_arr[1150] = 8'h0F;
		color_arr[1151] = 8'h0F;
		color_arr[1152] = 8'h0F;
		color_arr[1153] = 8'h0F;
		color_arr[1154] = 8'h0F;
		color_arr[1155] = 8'h0F;
		color_arr[1156] = 8'h0F;
		color_arr[1157] = 8'h0F;
		color_arr[1158] = 8'h0F;
		color_arr[1159] = 8'h0F;
		color_arr[1160] = 8'h0F;
		color_arr[1161] = 8'h0F;
		color_arr[1162] = 8'h0F;
		color_arr[1163] = 8'h0F;
		color_arr[1164] = 8'h0F;
		color_arr[1165] = 8'h0F;
		color_arr[1166] = 8'h0F;
		color_arr[1167] = 8'h0F;
		color_arr[1168] = 8'h0F;
		color_arr[1169] = 8'h0F;
		color_arr[1170] = 8'h0F;
		color_arr[1171] = 8'h0F;
		color_arr[1172] = 8'h0F;
		color_arr[1173] = 8'h0F;
		color_arr[1174] = 8'h0F;
		color_arr[1175] = 8'h0F;
		color_arr[1176] = 8'h0F;
		color_arr[1177] = 8'h0F;
		color_arr[1178] = 8'h0F;
		color_arr[1179] = 8'h0F;
		color_arr[1180] = 8'h0F;
		color_arr[1181] = 8'h0F;
		color_arr[1182] = 8'h0F;
		color_arr[1183] = 8'h0F;
		color_arr[1184] = 8'h0F;
		color_arr[1185] = 8'h0F;
		color_arr[1186] = 8'h0F;
		color_arr[1187] = 8'h0F;
		color_arr[1188] = 8'h0F;
		color_arr[1189] = 8'h0F;
		color_arr[1190] = 8'h0F;
		color_arr[1191] = 8'h0F;
		color_arr[1192] = 8'h0F;
		color_arr[1193] = 8'h0F;
		color_arr[1194] = 8'h0F;
		color_arr[1195] = 8'h0F;
		color_arr[1196] = 8'h0F;
		color_arr[1197] = 8'h0F;
		color_arr[1198] = 8'h0F;
		color_arr[1199] = 8'h0F;
		color_arr[1200] = 8'h0F;
		color_arr[1201] = 8'h0F;
		color_arr[1202] = 8'h0F;
		color_arr[1203] = 8'h0F;
		color_arr[1204] = 8'h0F;
		color_arr[1205] = 8'h0F;
		color_arr[1206] = 8'h0F;
		color_arr[1207] = 8'h0F;
		color_arr[1208] = 8'h0F;
		color_arr[1209] = 8'h0F;
		color_arr[1210] = 8'h0F;
		color_arr[1211] = 8'h0F;
		color_arr[1212] = 8'h0F;
		color_arr[1213] = 8'h0F;
		color_arr[1214] = 8'h0F;
		color_arr[1215] = 8'h0F;
		color_arr[1216] = 8'h0F;
		color_arr[1217] = 8'h0F;
		color_arr[1218] = 8'h0F;
		color_arr[1219] = 8'h0F;
		color_arr[1220] = 8'h0F;
		color_arr[1221] = 8'h0F;
		color_arr[1222] = 8'h0F;
		color_arr[1223] = 8'h0F;
		color_arr[1224] = 8'h0F;
		color_arr[1225] = 8'h0F;
		color_arr[1226] = 8'h0F;
		color_arr[1227] = 8'h0F;
		color_arr[1228] = 8'h0F;
		color_arr[1229] = 8'h0F;
		color_arr[1230] = 8'h0F;
		color_arr[1231] = 8'h0F;
		color_arr[1232] = 8'h0F;
		color_arr[1233] = 8'h0F;
		color_arr[1234] = 8'h0F;
		color_arr[1235] = 8'h0F;
		color_arr[1236] = 8'h0F;
		color_arr[1237] = 8'h0F;
		color_arr[1238] = 8'h0F;
		color_arr[1239] = 8'h0F;
		color_arr[1240] = 8'h0F;
		color_arr[1241] = 8'h0F;
		color_arr[1242] = 8'h0F;
		color_arr[1243] = 8'h0F;
		color_arr[1244] = 8'h0F;
		color_arr[1245] = 8'h0F;
		color_arr[1246] = 8'h0F;
		color_arr[1247] = 8'h0F;
		color_arr[1248] = 8'h0F;
		color_arr[1249] = 8'h0F;
		color_arr[1250] = 8'h0F;
		color_arr[1251] = 8'h0F;
		color_arr[1252] = 8'h0F;
		color_arr[1253] = 8'h0F;
		color_arr[1254] = 8'h0F;
		color_arr[1255] = 8'h0F;
		color_arr[1256] = 8'h0F;
		color_arr[1257] = 8'h0F;
		color_arr[1258] = 8'h0F;
		color_arr[1259] = 8'h0F;
		color_arr[1260] = 8'h0F;
		color_arr[1261] = 8'h0F;
		color_arr[1262] = 8'h0F;
		color_arr[1263] = 8'h0F;
		color_arr[1264] = 8'h0F;
		color_arr[1265] = 8'h0F;
		color_arr[1266] = 8'h0F;
		color_arr[1267] = 8'h0F;
		color_arr[1268] = 8'h0F;
		color_arr[1269] = 8'h0F;
		color_arr[1270] = 8'h0F;
		color_arr[1271] = 8'h0F;
		color_arr[1272] = 8'h0F;
		color_arr[1273] = 8'h0F;
		color_arr[1274] = 8'h0F;
		color_arr[1275] = 8'h0F;
		color_arr[1276] = 8'h0F;
		color_arr[1277] = 8'h0F;
		color_arr[1278] = 8'h0F;
		color_arr[1279] = 8'h0F;
		color_arr[1280] = 8'h0F;
		color_arr[1281] = 8'h0F;
		color_arr[1282] = 8'h0F;
		color_arr[1283] = 8'h0F;
		color_arr[1284] = 8'h0F;
		color_arr[1285] = 8'h0F;
		color_arr[1286] = 8'h0F;
		color_arr[1287] = 8'h0F;
		color_arr[1288] = 8'h0F;
		color_arr[1289] = 8'h0F;
		color_arr[1290] = 8'h0F;
		color_arr[1291] = 8'h0F;
		color_arr[1292] = 8'h0F;
		color_arr[1293] = 8'h0F;
		color_arr[1294] = 8'h0F;
		color_arr[1295] = 8'h0F;
		color_arr[1296] = 8'h0F;
		color_arr[1297] = 8'h0F;
		color_arr[1298] = 8'h0F;
		color_arr[1299] = 8'h0F;
		color_arr[1300] = 8'h0F;
		color_arr[1301] = 8'h0F;
		color_arr[1302] = 8'h0F;
		color_arr[1303] = 8'h0F;
		color_arr[1304] = 8'h0F;
		color_arr[1305] = 8'h0F;
		color_arr[1306] = 8'h0F;
		color_arr[1307] = 8'h0F;
		color_arr[1308] = 8'h0F;
		color_arr[1309] = 8'h0F;
		color_arr[1310] = 8'h0F;
		color_arr[1311] = 8'h0F;
		color_arr[1312] = 8'h0F;
		color_arr[1313] = 8'h0F;
		color_arr[1314] = 8'h0F;
		color_arr[1315] = 8'h0F;
		color_arr[1316] = 8'h0F;
		color_arr[1317] = 8'h0F;
		color_arr[1318] = 8'h0F;
		color_arr[1319] = 8'h0F;
		color_arr[1320] = 8'h0F;
		color_arr[1321] = 8'h0F;
		color_arr[1322] = 8'h0F;
		color_arr[1323] = 8'h0F;
		color_arr[1324] = 8'h0F;
		color_arr[1325] = 8'h0F;
		color_arr[1326] = 8'h0F;
		color_arr[1327] = 8'h0F;
		color_arr[1328] = 8'h0F;
		color_arr[1329] = 8'h0F;
		color_arr[1330] = 8'h0F;
		color_arr[1331] = 8'h0F;
		color_arr[1332] = 8'h0F;
		color_arr[1333] = 8'h0F;
		color_arr[1334] = 8'h0F;
		color_arr[1335] = 8'h0F;
		color_arr[1336] = 8'h0F;
		color_arr[1337] = 8'h0F;
		color_arr[1338] = 8'h0F;
		color_arr[1339] = 8'h0F;
		color_arr[1340] = 8'h0F;
		color_arr[1341] = 8'h0F;
		color_arr[1342] = 8'h0F;
		color_arr[1343] = 8'h0F;
		color_arr[1344] = 8'h0F;
		color_arr[1345] = 8'h0F;
		color_arr[1346] = 8'h0F;
		color_arr[1347] = 8'h0F;
		color_arr[1348] = 8'h0F;
		color_arr[1349] = 8'h0F;
		color_arr[1350] = 8'h0F;
		color_arr[1351] = 8'h0F;
		color_arr[1352] = 8'h0F;
		color_arr[1353] = 8'h0F;
		color_arr[1354] = 8'h0F;
		color_arr[1355] = 8'h0F;
		color_arr[1356] = 8'h0F;
		color_arr[1357] = 8'h0F;
		color_arr[1358] = 8'h0F;
		color_arr[1359] = 8'h0F;
		color_arr[1360] = 8'h0F;
		color_arr[1361] = 8'h0F;
		color_arr[1362] = 8'h0F;
		color_arr[1363] = 8'h0F;
		color_arr[1364] = 8'h0F;
		color_arr[1365] = 8'h0F;
		color_arr[1366] = 8'h0F;
		color_arr[1367] = 8'h0F;
		color_arr[1368] = 8'h0F;
		color_arr[1369] = 8'h0F;
		color_arr[1370] = 8'h0F;
		color_arr[1371] = 8'h0F;
		color_arr[1372] = 8'h0F;
		color_arr[1373] = 8'h0F;
		color_arr[1374] = 8'h0F;
		color_arr[1375] = 8'h0F;
		color_arr[1376] = 8'h0F;
		color_arr[1377] = 8'h0F;
		color_arr[1378] = 8'h0F;
		color_arr[1379] = 8'h0F;
		color_arr[1380] = 8'h0F;
		color_arr[1381] = 8'h0F;
		color_arr[1382] = 8'h0F;
		color_arr[1383] = 8'h0F;
		color_arr[1384] = 8'h0F;
		color_arr[1385] = 8'h0F;
		color_arr[1386] = 8'h0F;
		color_arr[1387] = 8'h0F;
		color_arr[1388] = 8'h0F;
		color_arr[1389] = 8'h0F;
		color_arr[1390] = 8'h0F;
		color_arr[1391] = 8'h0F;
		color_arr[1392] = 8'h0F;
		color_arr[1393] = 8'h0F;
		color_arr[1394] = 8'h0F;
		color_arr[1395] = 8'h0F;
		color_arr[1396] = 8'h0F;
		color_arr[1397] = 8'h0F;
		color_arr[1398] = 8'h0F;
		color_arr[1399] = 8'h0F;
		color_arr[1400] = 8'h0F;
		color_arr[1401] = 8'h0F;
		color_arr[1402] = 8'h0F;
		color_arr[1403] = 8'h0F;
		color_arr[1404] = 8'h0F;
		color_arr[1405] = 8'h0F;
		color_arr[1406] = 8'h0F;
		color_arr[1407] = 8'h0F;
		color_arr[1408] = 8'h0F;
		color_arr[1409] = 8'h0F;
		color_arr[1410] = 8'h0F;
		color_arr[1411] = 8'h0F;
		color_arr[1412] = 8'h0F;
		color_arr[1413] = 8'h0F;
		color_arr[1414] = 8'h0F;
		color_arr[1415] = 8'h0F;
		color_arr[1416] = 8'h0F;
		color_arr[1417] = 8'h0F;
		color_arr[1418] = 8'h0F;
		color_arr[1419] = 8'h0F;
		color_arr[1420] = 8'h0F;
		color_arr[1421] = 8'h0F;
		color_arr[1422] = 8'h0F;
		color_arr[1423] = 8'h0F;
		color_arr[1424] = 8'h0F;
		color_arr[1425] = 8'h0F;
		color_arr[1426] = 8'h0F;
		color_arr[1427] = 8'h0F;
		color_arr[1428] = 8'h0F;
		color_arr[1429] = 8'h0F;
		color_arr[1430] = 8'h0F;
		color_arr[1431] = 8'h0F;
		color_arr[1432] = 8'h0F;
		color_arr[1433] = 8'h0F;
		color_arr[1434] = 8'h0F;
		color_arr[1435] = 8'h0F;
		color_arr[1436] = 8'h0F;
		color_arr[1437] = 8'h0F;
		color_arr[1438] = 8'h0F;
		color_arr[1439] = 8'h0F;
		color_arr[1440] = 8'h0F;
		color_arr[1441] = 8'h0F;
		color_arr[1442] = 8'h0F;
		color_arr[1443] = 8'h0F;
		color_arr[1444] = 8'h0F;
		color_arr[1445] = 8'h0F;
		color_arr[1446] = 8'h0F;
		color_arr[1447] = 8'h0F;
		color_arr[1448] = 8'h0F;
		color_arr[1449] = 8'h0F;
		color_arr[1450] = 8'h0F;
		color_arr[1451] = 8'h0F;
		color_arr[1452] = 8'h0F;
		color_arr[1453] = 8'h0F;
		color_arr[1454] = 8'h0F;
		color_arr[1455] = 8'h0F;
		color_arr[1456] = 8'h0F;
		color_arr[1457] = 8'h0F;
		color_arr[1458] = 8'h0F;
		color_arr[1459] = 8'h0F;
		color_arr[1460] = 8'h0F;
		color_arr[1461] = 8'h0F;
		color_arr[1462] = 8'h0F;
		color_arr[1463] = 8'h0F;
		color_arr[1464] = 8'h0F;
		color_arr[1465] = 8'h0F;
		color_arr[1466] = 8'h0F;
		color_arr[1467] = 8'h0F;
		color_arr[1468] = 8'h0F;
		color_arr[1469] = 8'h0F;
		color_arr[1470] = 8'h0F;
		color_arr[1471] = 8'h0F;
		color_arr[1472] = 8'h0F;
		color_arr[1473] = 8'h0F;
		color_arr[1474] = 8'h0F;
		color_arr[1475] = 8'h0F;
		color_arr[1476] = 8'h0F;
		color_arr[1477] = 8'h0F;
		color_arr[1478] = 8'h0F;
		color_arr[1479] = 8'h0F;
		color_arr[1480] = 8'h0F;
		color_arr[1481] = 8'h0F;
		color_arr[1482] = 8'h0F;
		color_arr[1483] = 8'h0F;
		color_arr[1484] = 8'h0F;
		color_arr[1485] = 8'h0F;
		color_arr[1486] = 8'h0F;
		color_arr[1487] = 8'h0F;
		color_arr[1488] = 8'h0F;
		color_arr[1489] = 8'h0F;
		color_arr[1490] = 8'h0F;
		color_arr[1491] = 8'h0F;
		color_arr[1492] = 8'h0F;
		color_arr[1493] = 8'h0F;
		color_arr[1494] = 8'h0F;
		color_arr[1495] = 8'h0F;
		color_arr[1496] = 8'h0F;
		color_arr[1497] = 8'h0F;
		color_arr[1498] = 8'h0F;
		color_arr[1499] = 8'h0F;
		color_arr[1500] = 8'h0F;
		color_arr[1501] = 8'h0F;
		color_arr[1502] = 8'h0F;
		color_arr[1503] = 8'h0F;
		color_arr[1504] = 8'h0F;
		color_arr[1505] = 8'h0F;
		color_arr[1506] = 8'h0F;
		color_arr[1507] = 8'h0F;
		color_arr[1508] = 8'h0F;
		color_arr[1509] = 8'h0F;
		color_arr[1510] = 8'h0F;
		color_arr[1511] = 8'h0F;
		color_arr[1512] = 8'h0F;
		color_arr[1513] = 8'h0F;
		color_arr[1514] = 8'h0F;
		color_arr[1515] = 8'h0F;
		color_arr[1516] = 8'h0F;
		color_arr[1517] = 8'h0F;
		color_arr[1518] = 8'h0F;
		color_arr[1519] = 8'h0F;
		color_arr[1520] = 8'h0F;
		color_arr[1521] = 8'h0F;
		color_arr[1522] = 8'h0F;
		color_arr[1523] = 8'h0F;
		color_arr[1524] = 8'h0F;
		color_arr[1525] = 8'h0F;
		color_arr[1526] = 8'h0F;
		color_arr[1527] = 8'h0F;
		color_arr[1528] = 8'h0F;
		color_arr[1529] = 8'h0F;
		color_arr[1530] = 8'h0F;
		color_arr[1531] = 8'h0F;
		color_arr[1532] = 8'h0F;
		color_arr[1533] = 8'h0F;
		color_arr[1534] = 8'h0F;
		color_arr[1535] = 8'h0F;
		color_arr[1536] = 8'h0F;
		color_arr[1537] = 8'h0F;
		color_arr[1538] = 8'h0F;
		color_arr[1539] = 8'h0F;
		color_arr[1540] = 8'h0F;
		color_arr[1541] = 8'h0F;
		color_arr[1542] = 8'h0F;
		color_arr[1543] = 8'h0F;
		color_arr[1544] = 8'h0F;
		color_arr[1545] = 8'h0F;
		color_arr[1546] = 8'h0F;
		color_arr[1547] = 8'h0F;
		color_arr[1548] = 8'h0F;
		color_arr[1549] = 8'h0F;
		color_arr[1550] = 8'h0F;
		color_arr[1551] = 8'h0F;
		color_arr[1552] = 8'h0F;
		color_arr[1553] = 8'h0F;
		color_arr[1554] = 8'h0F;
		color_arr[1555] = 8'h0F;
		color_arr[1556] = 8'h0F;
		color_arr[1557] = 8'h0F;
		color_arr[1558] = 8'h0F;
		color_arr[1559] = 8'h0F;
		color_arr[1560] = 8'h0F;
		color_arr[1561] = 8'h0F;
		color_arr[1562] = 8'h0F;
		color_arr[1563] = 8'h0F;
		color_arr[1564] = 8'h0F;
		color_arr[1565] = 8'h0F;
		color_arr[1566] = 8'h0F;
		color_arr[1567] = 8'h0F;
		color_arr[1568] = 8'h0F;
		color_arr[1569] = 8'h0F;
		color_arr[1570] = 8'h0F;
		color_arr[1571] = 8'h0F;
		color_arr[1572] = 8'h0F;
		color_arr[1573] = 8'h0F;
		color_arr[1574] = 8'h0F;
		color_arr[1575] = 8'h0F;
		color_arr[1576] = 8'h0F;
		color_arr[1577] = 8'h0F;
		color_arr[1578] = 8'h0F;
		color_arr[1579] = 8'h0F;
		color_arr[1580] = 8'h0F;
		color_arr[1581] = 8'h0F;
		color_arr[1582] = 8'h0F;
		color_arr[1583] = 8'h0F;
		color_arr[1584] = 8'h0F;
		color_arr[1585] = 8'h0F;
		color_arr[1586] = 8'h0F;
		color_arr[1587] = 8'h0F;
		color_arr[1588] = 8'h0F;
		color_arr[1589] = 8'h0F;
		color_arr[1590] = 8'h0F;
		color_arr[1591] = 8'h0F;
		color_arr[1592] = 8'h0F;
		color_arr[1593] = 8'h0F;
		color_arr[1594] = 8'h0F;
		color_arr[1595] = 8'h0F;
		color_arr[1596] = 8'h0F;
		color_arr[1597] = 8'h0F;
		color_arr[1598] = 8'h0F;
		color_arr[1599] = 8'h0F;
		color_arr[1600] = 8'h0F;
		color_arr[1601] = 8'h0F;
		color_arr[1602] = 8'h0F;
		color_arr[1603] = 8'h0F;
		color_arr[1604] = 8'h0F;
		color_arr[1605] = 8'h0F;
		color_arr[1606] = 8'h0F;
		color_arr[1607] = 8'h0F;
		color_arr[1608] = 8'h0F;
		color_arr[1609] = 8'h0F;
		color_arr[1610] = 8'h0F;
		color_arr[1611] = 8'h0F;
		color_arr[1612] = 8'h0F;
		color_arr[1613] = 8'h0F;
		color_arr[1614] = 8'h0F;
		color_arr[1615] = 8'h0F;
		color_arr[1616] = 8'h0F;
		color_arr[1617] = 8'h0F;
		color_arr[1618] = 8'h0F;
		color_arr[1619] = 8'h0F;
		color_arr[1620] = 8'h0F;
		color_arr[1621] = 8'h0F;
		color_arr[1622] = 8'h0F;
		color_arr[1623] = 8'h0F;
		color_arr[1624] = 8'h0F;
		color_arr[1625] = 8'h0F;
		color_arr[1626] = 8'h0F;
		color_arr[1627] = 8'h0F;
		color_arr[1628] = 8'h0F;
		color_arr[1629] = 8'h0F;
		color_arr[1630] = 8'h0F;
		color_arr[1631] = 8'h0F;
		color_arr[1632] = 8'h0F;
		color_arr[1633] = 8'h0F;
		color_arr[1634] = 8'h0F;
		color_arr[1635] = 8'h0F;
		color_arr[1636] = 8'h0F;
		color_arr[1637] = 8'h0F;
		color_arr[1638] = 8'h0F;
		color_arr[1639] = 8'h0F;
		color_arr[1640] = 8'h0F;
		color_arr[1641] = 8'h0F;
		color_arr[1642] = 8'h0F;
		color_arr[1643] = 8'h0F;
		color_arr[1644] = 8'h0F;
		color_arr[1645] = 8'h0F;
		color_arr[1646] = 8'h0F;
		color_arr[1647] = 8'h0F;
		color_arr[1648] = 8'h0F;
		color_arr[1649] = 8'h0F;
		color_arr[1650] = 8'h0F;
		color_arr[1651] = 8'h0F;
		color_arr[1652] = 8'h0F;
		color_arr[1653] = 8'h0F;
		color_arr[1654] = 8'h0F;
		color_arr[1655] = 8'h0F;
		color_arr[1656] = 8'h0F;
		color_arr[1657] = 8'h0F;
		color_arr[1658] = 8'h0F;
		color_arr[1659] = 8'h0F;
		color_arr[1660] = 8'h0F;
		color_arr[1661] = 8'h0F;
		color_arr[1662] = 8'h0F;
		color_arr[1663] = 8'h0F;
		color_arr[1664] = 8'h0F;
		color_arr[1665] = 8'h0F;
		color_arr[1666] = 8'h0F;
		color_arr[1667] = 8'h0F;
		color_arr[1668] = 8'h0F;
		color_arr[1669] = 8'h0F;
		color_arr[1670] = 8'h0F;
		color_arr[1671] = 8'h0F;
		color_arr[1672] = 8'h0F;
		color_arr[1673] = 8'h0F;
		color_arr[1674] = 8'h0F;
		color_arr[1675] = 8'h0F;
		color_arr[1676] = 8'h0F;
		color_arr[1677] = 8'h0F;
		color_arr[1678] = 8'h0F;
		color_arr[1679] = 8'h0F;
		color_arr[1680] = 8'h0F;
		color_arr[1681] = 8'h0F;
		color_arr[1682] = 8'h0F;
		color_arr[1683] = 8'h0F;
		color_arr[1684] = 8'h0F;
		color_arr[1685] = 8'h0F;
		color_arr[1686] = 8'h0F;
		color_arr[1687] = 8'h0F;
		color_arr[1688] = 8'h0F;
		color_arr[1689] = 8'h0F;
		color_arr[1690] = 8'h0F;
		color_arr[1691] = 8'h0F;
		color_arr[1692] = 8'h0F;
		color_arr[1693] = 8'h0F;
		color_arr[1694] = 8'h0F;
		color_arr[1695] = 8'h0F;
		color_arr[1696] = 8'h0F;
		color_arr[1697] = 8'h0F;
		color_arr[1698] = 8'h0F;
		color_arr[1699] = 8'h0F;
		color_arr[1700] = 8'h0F;
		color_arr[1701] = 8'h0F;
		color_arr[1702] = 8'h0F;
		color_arr[1703] = 8'h0F;
		color_arr[1704] = 8'h0F;
		color_arr[1705] = 8'h0F;
		color_arr[1706] = 8'h0F;
		color_arr[1707] = 8'h0F;
		color_arr[1708] = 8'h0F;
		color_arr[1709] = 8'h0F;
		color_arr[1710] = 8'h0F;
		color_arr[1711] = 8'h0F;
		color_arr[1712] = 8'h0F;
		color_arr[1713] = 8'h0F;
		color_arr[1714] = 8'h0F;
		color_arr[1715] = 8'h0F;
		color_arr[1716] = 8'h0F;
		color_arr[1717] = 8'h0F;
		color_arr[1718] = 8'h0F;
		color_arr[1719] = 8'h0F;
		color_arr[1720] = 8'h0F;
		color_arr[1721] = 8'h0F;
		color_arr[1722] = 8'h0F;
		color_arr[1723] = 8'h0F;
		color_arr[1724] = 8'h0F;
		color_arr[1725] = 8'h0F;
		color_arr[1726] = 8'h0F;
		color_arr[1727] = 8'h0F;
		color_arr[1728] = 8'h0F;
		color_arr[1729] = 8'h0F;
		color_arr[1730] = 8'h0F;
		color_arr[1731] = 8'h0F;
		color_arr[1732] = 8'h0F;
		color_arr[1733] = 8'h0F;
		color_arr[1734] = 8'h0F;
		color_arr[1735] = 8'h0F;
		color_arr[1736] = 8'h0F;
		color_arr[1737] = 8'h0F;
		color_arr[1738] = 8'h0F;
		color_arr[1739] = 8'h0F;
		color_arr[1740] = 8'h0F;
		color_arr[1741] = 8'h0F;
		color_arr[1742] = 8'h0F;
		color_arr[1743] = 8'h0F;
		color_arr[1744] = 8'h0F;
		color_arr[1745] = 8'h0F;
		color_arr[1746] = 8'h0F;
		color_arr[1747] = 8'h0F;
		color_arr[1748] = 8'h0F;
		color_arr[1749] = 8'h0F;
		color_arr[1750] = 8'h0F;
		color_arr[1751] = 8'h0F;
		color_arr[1752] = 8'h0F;
		color_arr[1753] = 8'h0F;
		color_arr[1754] = 8'h0F;
		color_arr[1755] = 8'h0F;
		color_arr[1756] = 8'h0F;
		color_arr[1757] = 8'h0F;
		color_arr[1758] = 8'h0F;
		color_arr[1759] = 8'h0F;
		color_arr[1760] = 8'h0F;
		color_arr[1761] = 8'h0F;
		color_arr[1762] = 8'h0F;
		color_arr[1763] = 8'h0F;
		color_arr[1764] = 8'h0F;
		color_arr[1765] = 8'h0F;
		color_arr[1766] = 8'h0F;
		color_arr[1767] = 8'h0F;
		color_arr[1768] = 8'h0F;
		color_arr[1769] = 8'h0F;
		color_arr[1770] = 8'h0F;
		color_arr[1771] = 8'h0F;
		color_arr[1772] = 8'h0F;
		color_arr[1773] = 8'h0F;
		color_arr[1774] = 8'h0F;
		color_arr[1775] = 8'h0F;
		color_arr[1776] = 8'h0F;
		color_arr[1777] = 8'h0F;
		color_arr[1778] = 8'h0F;
		color_arr[1779] = 8'h0F;
		color_arr[1780] = 8'h0F;
		color_arr[1781] = 8'h0F;
		color_arr[1782] = 8'h0F;
		color_arr[1783] = 8'h0F;
		color_arr[1784] = 8'h0F;
		color_arr[1785] = 8'h0F;
		color_arr[1786] = 8'h0F;
		color_arr[1787] = 8'h0F;
		color_arr[1788] = 8'h0F;
		color_arr[1789] = 8'h0F;
		color_arr[1790] = 8'h0F;
		color_arr[1791] = 8'h0F;
		color_arr[1792] = 8'h0F;
		color_arr[1793] = 8'h0F;
		color_arr[1794] = 8'h0F;
		color_arr[1795] = 8'h0F;
		color_arr[1796] = 8'h0F;
		color_arr[1797] = 8'h0F;
		color_arr[1798] = 8'h0F;
		color_arr[1799] = 8'h0F;
		color_arr[1800] = 8'h0F;
		color_arr[1801] = 8'h0F;
		color_arr[1802] = 8'h0F;
		color_arr[1803] = 8'h0F;
		color_arr[1804] = 8'h0F;
		color_arr[1805] = 8'h0F;
		color_arr[1806] = 8'h0F;
		color_arr[1807] = 8'h0F;
		color_arr[1808] = 8'h0F;
		color_arr[1809] = 8'h0F;
		color_arr[1810] = 8'h0F;
		color_arr[1811] = 8'h0F;
		color_arr[1812] = 8'h0F;
		color_arr[1813] = 8'h0F;
		color_arr[1814] = 8'h0F;
		color_arr[1815] = 8'h0F;
		color_arr[1816] = 8'h0F;
		color_arr[1817] = 8'h0F;
		color_arr[1818] = 8'h0F;
		color_arr[1819] = 8'h0F;
		color_arr[1820] = 8'h0F;
		color_arr[1821] = 8'h0F;
		color_arr[1822] = 8'h0F;
		color_arr[1823] = 8'h0F;
		color_arr[1824] = 8'h0F;
		color_arr[1825] = 8'h0F;
		color_arr[1826] = 8'h0F;
		color_arr[1827] = 8'h0F;
		color_arr[1828] = 8'h0F;
		color_arr[1829] = 8'h0F;
		color_arr[1830] = 8'h0F;
		color_arr[1831] = 8'h0F;
		color_arr[1832] = 8'h0F;
		color_arr[1833] = 8'h0F;
		color_arr[1834] = 8'h0F;
		color_arr[1835] = 8'h0F;
		color_arr[1836] = 8'h0F;
		color_arr[1837] = 8'h0F;
		color_arr[1838] = 8'h0F;
		color_arr[1839] = 8'h0F;
		color_arr[1840] = 8'h0F;
		color_arr[1841] = 8'h0F;
		color_arr[1842] = 8'h0F;
		color_arr[1843] = 8'h0F;
		color_arr[1844] = 8'h0F;
		color_arr[1845] = 8'h0F;
		color_arr[1846] = 8'h0F;
		color_arr[1847] = 8'h0F;
		color_arr[1848] = 8'h0F;
		color_arr[1849] = 8'h0F;
		color_arr[1850] = 8'h0F;
		color_arr[1851] = 8'h0F;
		color_arr[1852] = 8'h0F;
		color_arr[1853] = 8'h0F;
		color_arr[1854] = 8'h0F;
		color_arr[1855] = 8'h0F;
		color_arr[1856] = 8'h0F;
		color_arr[1857] = 8'h0F;
		color_arr[1858] = 8'h0F;
		color_arr[1859] = 8'h0F;
		color_arr[1860] = 8'h0F;
		color_arr[1861] = 8'h0F;
		color_arr[1862] = 8'h0F;
		color_arr[1863] = 8'h0F;
		color_arr[1864] = 8'h0F;
		color_arr[1865] = 8'h0F;
		color_arr[1866] = 8'h0F;
		color_arr[1867] = 8'h0F;
		color_arr[1868] = 8'h0F;
		color_arr[1869] = 8'h0F;
		color_arr[1870] = 8'h0F;
		color_arr[1871] = 8'h0F;
		color_arr[1872] = 8'h0F;
		color_arr[1873] = 8'h0F;
		color_arr[1874] = 8'h0F;
		color_arr[1875] = 8'h0F;
		color_arr[1876] = 8'h0F;
		color_arr[1877] = 8'h0F;
		color_arr[1878] = 8'h0F;
		color_arr[1879] = 8'h0F;
		color_arr[1880] = 8'h0F;
		color_arr[1881] = 8'h0F;
		color_arr[1882] = 8'h0F;
		color_arr[1883] = 8'h0F;
		color_arr[1884] = 8'h0F;
		color_arr[1885] = 8'h0F;
		color_arr[1886] = 8'h0F;
		color_arr[1887] = 8'h0F;
		color_arr[1888] = 8'h0F;
		color_arr[1889] = 8'h0F;
		color_arr[1890] = 8'h0F;
		color_arr[1891] = 8'h0F;
		color_arr[1892] = 8'h0F;
		color_arr[1893] = 8'h0F;
		color_arr[1894] = 8'h0F;
		color_arr[1895] = 8'h0F;
		color_arr[1896] = 8'h0F;
		color_arr[1897] = 8'h0F;
		color_arr[1898] = 8'h0F;
		color_arr[1899] = 8'h0F;
		color_arr[1900] = 8'h0F;
		color_arr[1901] = 8'h0F;
		color_arr[1902] = 8'h0F;
		color_arr[1903] = 8'h0F;
		color_arr[1904] = 8'h0F;
		color_arr[1905] = 8'h0F;
		color_arr[1906] = 8'h0F;
		color_arr[1907] = 8'h0F;
		color_arr[1908] = 8'h0F;
		color_arr[1909] = 8'h0F;
		color_arr[1910] = 8'h0F;
		color_arr[1911] = 8'h0F;
		color_arr[1912] = 8'h0F;
		color_arr[1913] = 8'h0F;
		color_arr[1914] = 8'h0F;
		color_arr[1915] = 8'h0F;
		color_arr[1916] = 8'h0F;
		color_arr[1917] = 8'h0F;
		color_arr[1918] = 8'h0F;
		color_arr[1919] = 8'h0F;
		color_arr[1920] = 8'h0F;
		color_arr[1921] = 8'h0F;
		color_arr[1922] = 8'h0F;
		color_arr[1923] = 8'h0F;
		color_arr[1924] = 8'h0F;
		color_arr[1925] = 8'h0F;
		color_arr[1926] = 8'h0F;
		color_arr[1927] = 8'h0F;
		color_arr[1928] = 8'h0F;
		color_arr[1929] = 8'h0F;
		color_arr[1930] = 8'h0F;
		color_arr[1931] = 8'h0F;
		color_arr[1932] = 8'h0F;
		color_arr[1933] = 8'h0F;
		color_arr[1934] = 8'h0F;
		color_arr[1935] = 8'h0F;
		color_arr[1936] = 8'h0F;
		color_arr[1937] = 8'h0F;
		color_arr[1938] = 8'h0F;
		color_arr[1939] = 8'h0F;
		color_arr[1940] = 8'h0F;
		color_arr[1941] = 8'h0F;
		color_arr[1942] = 8'h0F;
		color_arr[1943] = 8'h0F;
		color_arr[1944] = 8'h0F;
		color_arr[1945] = 8'h0F;
		color_arr[1946] = 8'h0F;
		color_arr[1947] = 8'h0F;
		color_arr[1948] = 8'h0F;
		color_arr[1949] = 8'h0F;
		color_arr[1950] = 8'h0F;
		color_arr[1951] = 8'h0F;
		color_arr[1952] = 8'h0F;
		color_arr[1953] = 8'h0F;
		color_arr[1954] = 8'h0F;
		color_arr[1955] = 8'h0F;
		color_arr[1956] = 8'h0F;
		color_arr[1957] = 8'h0F;
		color_arr[1958] = 8'h0F;
		color_arr[1959] = 8'h0F;
		color_arr[1960] = 8'h0F;
		color_arr[1961] = 8'h0F;
		color_arr[1962] = 8'h0F;
		color_arr[1963] = 8'h0F;
		color_arr[1964] = 8'h0F;
		color_arr[1965] = 8'h0F;
		color_arr[1966] = 8'h0F;
		color_arr[1967] = 8'h0F;
		color_arr[1968] = 8'h0F;
		color_arr[1969] = 8'h0F;
		color_arr[1970] = 8'h0F;
		color_arr[1971] = 8'h0F;
		color_arr[1972] = 8'h0F;
		color_arr[1973] = 8'h0F;
		color_arr[1974] = 8'h0F;
		color_arr[1975] = 8'h0F;
		color_arr[1976] = 8'h0F;
		color_arr[1977] = 8'h0F;
		color_arr[1978] = 8'h0F;
		color_arr[1979] = 8'h0F;
		color_arr[1980] = 8'h0F;
		color_arr[1981] = 8'h0F;
		color_arr[1982] = 8'h0F;
		color_arr[1983] = 8'h0F;
		color_arr[1984] = 8'h0F;
		color_arr[1985] = 8'h0F;
		color_arr[1986] = 8'h0F;
		color_arr[1987] = 8'h0F;
		color_arr[1988] = 8'h0F;
		color_arr[1989] = 8'h0F;
		color_arr[1990] = 8'h0F;
		color_arr[1991] = 8'h0F;
		color_arr[1992] = 8'h0F;
		color_arr[1993] = 8'h0F;
		color_arr[1994] = 8'h0F;
		color_arr[1995] = 8'h0F;
		color_arr[1996] = 8'h0F;
		color_arr[1997] = 8'h0F;
		color_arr[1998] = 8'h0F;
		color_arr[1999] = 8'h0F;
		color_arr[2000] = 8'h0F;
		color_arr[2001] = 8'h0F;
		color_arr[2002] = 8'h0F;
		color_arr[2003] = 8'h0F;
		color_arr[2004] = 8'h0F;
		color_arr[2005] = 8'h0F;
		color_arr[2006] = 8'h0F;
		color_arr[2007] = 8'h0F;
		color_arr[2008] = 8'h0F;
		color_arr[2009] = 8'h0F;
		color_arr[2010] = 8'h0F;
		color_arr[2011] = 8'h0F;
		color_arr[2012] = 8'h0F;
		color_arr[2013] = 8'h0F;
		color_arr[2014] = 8'h0F;
		color_arr[2015] = 8'h0F;
		color_arr[2016] = 8'h0F;
		color_arr[2017] = 8'h0F;
		color_arr[2018] = 8'h0F;
		color_arr[2019] = 8'h0F;
		color_arr[2020] = 8'h0F;
		color_arr[2021] = 8'h0F;
		color_arr[2022] = 8'h0F;
		color_arr[2023] = 8'h0F;
		color_arr[2024] = 8'h0F;
		color_arr[2025] = 8'h0F;
		color_arr[2026] = 8'h0F;
		color_arr[2027] = 8'h0F;
		color_arr[2028] = 8'h0F;
		color_arr[2029] = 8'h0F;
		color_arr[2030] = 8'h0F;
		color_arr[2031] = 8'h0F;
		color_arr[2032] = 8'h0F;
		color_arr[2033] = 8'h0F;
		color_arr[2034] = 8'h0F;
		color_arr[2035] = 8'h0F;
		color_arr[2036] = 8'h0F;
		color_arr[2037] = 8'h0F;
		color_arr[2038] = 8'h0F;
		color_arr[2039] = 8'h0F;
		color_arr[2040] = 8'h0F;
		color_arr[2041] = 8'h0F;
		color_arr[2042] = 8'h0F;
		color_arr[2043] = 8'h0F;
		color_arr[2044] = 8'h0F;
		color_arr[2045] = 8'h0F;
		color_arr[2046] = 8'h0F;
		color_arr[2047] = 8'h0F;
	end

	always @(posedge clk) begin
		color_out <= color_arr[addr][5:0];
	end
endmodule
