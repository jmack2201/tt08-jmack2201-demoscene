module pwm (
    input clk, rst_n, audio_in,
    output pwm_out
);
    
endmodule