module audio_source (
    input clk, rst_n,
    input [1:0] audio_select,
    output audio_out
);
    
endmodule