module sprite_rom0 (
	input clk,
	input [11:0] addr,
	output reg [5:0] color_out
);
	reg [5:0] color_arr [SPRITE_SIZE*SPRITE_SIZE-1:0];

	initial begin
		color_arr[0] = 8'b00010010;
		color_arr[1] = 8'b00010010;
		color_arr[2] = 8'b00010010;
		color_arr[3] = 8'b00010010;
		color_arr[4] = 8'b00010010;
		color_arr[5] = 8'b00010010;
		color_arr[6] = 8'b00010010;
		color_arr[7] = 8'b00010010;
		color_arr[8] = 8'b00010010;
		color_arr[9] = 8'b00010010;
		color_arr[10] = 8'b00010010;
		color_arr[11] = 8'b00010010;
		color_arr[12] = 8'b00010010;
		color_arr[13] = 8'b00010010;
		color_arr[14] = 8'b00010010;
		color_arr[15] = 8'b00010010;
		color_arr[16] = 8'b00010010;
		color_arr[17] = 8'b00010010;
		color_arr[18] = 8'b00010010;
		color_arr[19] = 8'b00010010;
		color_arr[20] = 8'b00010010;
		color_arr[21] = 8'b00010010;
		color_arr[22] = 8'b00010010;
		color_arr[23] = 8'b00010010;
		color_arr[24] = 8'b00010010;
		color_arr[25] = 8'b00010010;
		color_arr[26] = 8'b00010010;
		color_arr[27] = 8'b00010010;
		color_arr[28] = 8'b00010010;
		color_arr[29] = 8'b00010010;
		color_arr[30] = 8'b00010010;
		color_arr[31] = 8'b00010010;
		color_arr[32] = 8'b00010010;
		color_arr[33] = 8'b00010010;
		color_arr[34] = 8'b00010010;
		color_arr[35] = 8'b00010010;
		color_arr[36] = 8'b00010010;
		color_arr[37] = 8'b00010010;
		color_arr[38] = 8'b00010010;
		color_arr[39] = 8'b00010010;
		color_arr[40] = 8'b00010010;
		color_arr[41] = 8'b00010010;
		color_arr[42] = 8'b00010010;
		color_arr[43] = 8'b00010010;
		color_arr[44] = 8'b00010010;
		color_arr[45] = 8'b00010010;
		color_arr[46] = 8'b00010010;
		color_arr[47] = 8'b00010010;
		color_arr[48] = 8'b00010010;
		color_arr[49] = 8'b00010010;
		color_arr[50] = 8'b00010010;
		color_arr[51] = 8'b00010010;
		color_arr[52] = 8'b00010010;
		color_arr[53] = 8'b00010010;
		color_arr[54] = 8'b00010010;
		color_arr[55] = 8'b00010010;
		color_arr[56] = 8'b00010010;
		color_arr[57] = 8'b00010010;
		color_arr[58] = 8'b00010010;
		color_arr[59] = 8'b00010010;
		color_arr[60] = 8'b00010010;
		color_arr[61] = 8'b00010010;
		color_arr[62] = 8'b00010010;
		color_arr[63] = 8'b00010010;
		color_arr[64] = 8'b00010010;
		color_arr[65] = 8'b00010010;
		color_arr[66] = 8'b00010010;
		color_arr[67] = 8'b00010010;
		color_arr[68] = 8'b00010010;
		color_arr[69] = 8'b00010010;
		color_arr[70] = 8'b00010010;
		color_arr[71] = 8'b00010010;
		color_arr[72] = 8'b00010010;
		color_arr[73] = 8'b00010010;
		color_arr[74] = 8'b00010010;
		color_arr[75] = 8'b00010010;
		color_arr[76] = 8'b00010010;
		color_arr[77] = 8'b00010010;
		color_arr[78] = 8'b00010010;
		color_arr[79] = 8'b00010010;
		color_arr[80] = 8'b00010010;
		color_arr[81] = 8'b00010010;
		color_arr[82] = 8'b00010010;
		color_arr[83] = 8'b00010010;
		color_arr[84] = 8'b00010010;
		color_arr[85] = 8'b00010010;
		color_arr[86] = 8'b00010010;
		color_arr[87] = 8'b00010010;
		color_arr[88] = 8'b00010010;
		color_arr[89] = 8'b00010010;
		color_arr[90] = 8'b00010010;
		color_arr[91] = 8'b00010010;
		color_arr[92] = 8'b00010010;
		color_arr[93] = 8'b00010010;
		color_arr[94] = 8'b00010010;
		color_arr[95] = 8'b00010010;
		color_arr[96] = 8'b00010010;
		color_arr[97] = 8'b00010010;
		color_arr[98] = 8'b00010010;
		color_arr[99] = 8'b00010010;
		color_arr[100] = 8'b00010010;
		color_arr[101] = 8'b00010010;
		color_arr[102] = 8'b00010010;
		color_arr[103] = 8'b00010010;
		color_arr[104] = 8'b00010010;
		color_arr[105] = 8'b00010010;
		color_arr[106] = 8'b00010010;
		color_arr[107] = 8'b00010010;
		color_arr[108] = 8'b00010010;
		color_arr[109] = 8'b00010010;
		color_arr[110] = 8'b00010010;
		color_arr[111] = 8'b00010010;
		color_arr[112] = 8'b00010010;
		color_arr[113] = 8'b00010010;
		color_arr[114] = 8'b00010010;
		color_arr[115] = 8'b00010010;
		color_arr[116] = 8'b00010010;
		color_arr[117] = 8'b00010010;
		color_arr[118] = 8'b00010010;
		color_arr[119] = 8'b00010010;
		color_arr[120] = 8'b00010010;
		color_arr[121] = 8'b00010010;
		color_arr[122] = 8'b00010010;
		color_arr[123] = 8'b00000000;
		color_arr[124] = 8'b00000000;
		color_arr[125] = 8'b00000000;
		color_arr[126] = 8'b00000000;
		color_arr[127] = 8'b00000000;
		color_arr[128] = 8'b00010010;
		color_arr[129] = 8'b00010010;
		color_arr[130] = 8'b00010010;
		color_arr[131] = 8'b00010010;
		color_arr[132] = 8'b00010010;
		color_arr[133] = 8'b00010010;
		color_arr[134] = 8'b00010010;
		color_arr[135] = 8'b00010010;
		color_arr[136] = 8'b00010010;
		color_arr[137] = 8'b00010010;
		color_arr[138] = 8'b00010010;
		color_arr[139] = 8'b00010010;
		color_arr[140] = 8'b00010010;
		color_arr[141] = 8'b00010010;
		color_arr[142] = 8'b00010010;
		color_arr[143] = 8'b00010010;
		color_arr[144] = 8'b00010010;
		color_arr[145] = 8'b00010010;
		color_arr[146] = 8'b00010010;
		color_arr[147] = 8'b00010010;
		color_arr[148] = 8'b00010010;
		color_arr[149] = 8'b00010010;
		color_arr[150] = 8'b00010010;
		color_arr[151] = 8'b00010010;
		color_arr[152] = 8'b00010010;
		color_arr[153] = 8'b00010010;
		color_arr[154] = 8'b00010010;
		color_arr[155] = 8'b00010010;
		color_arr[156] = 8'b00010010;
		color_arr[157] = 8'b00010010;
		color_arr[158] = 8'b00010010;
		color_arr[159] = 8'b00010010;
		color_arr[160] = 8'b00010010;
		color_arr[161] = 8'b00010010;
		color_arr[162] = 8'b00010010;
		color_arr[163] = 8'b00010010;
		color_arr[164] = 8'b00010010;
		color_arr[165] = 8'b00010010;
		color_arr[166] = 8'b00010010;
		color_arr[167] = 8'b00010010;
		color_arr[168] = 8'b00010010;
		color_arr[169] = 8'b00010010;
		color_arr[170] = 8'b00010010;
		color_arr[171] = 8'b00010010;
		color_arr[172] = 8'b00010010;
		color_arr[173] = 8'b00010010;
		color_arr[174] = 8'b00010010;
		color_arr[175] = 8'b00010010;
		color_arr[176] = 8'b00010010;
		color_arr[177] = 8'b00010010;
		color_arr[178] = 8'b00010010;
		color_arr[179] = 8'b00010010;
		color_arr[180] = 8'b00010010;
		color_arr[181] = 8'b00010010;
		color_arr[182] = 8'b00010010;
		color_arr[183] = 8'b00010010;
		color_arr[184] = 8'b00000000;
		color_arr[185] = 8'b00000000;
		color_arr[186] = 8'b00000000;
		color_arr[187] = 8'b00000000;
		color_arr[188] = 8'b00000000;
		color_arr[189] = 8'b00000000;
		color_arr[190] = 8'b00000000;
		color_arr[191] = 8'b00000000;
		color_arr[192] = 8'b00010010;
		color_arr[193] = 8'b00010010;
		color_arr[194] = 8'b00010010;
		color_arr[195] = 8'b00010010;
		color_arr[196] = 8'b00010010;
		color_arr[197] = 8'b00010010;
		color_arr[198] = 8'b00010010;
		color_arr[199] = 8'b00010010;
		color_arr[200] = 8'b00010010;
		color_arr[201] = 8'b00010010;
		color_arr[202] = 8'b00010010;
		color_arr[203] = 8'b00010010;
		color_arr[204] = 8'b00010010;
		color_arr[205] = 8'b00010010;
		color_arr[206] = 8'b00010010;
		color_arr[207] = 8'b00010010;
		color_arr[208] = 8'b00010010;
		color_arr[209] = 8'b00010010;
		color_arr[210] = 8'b00010010;
		color_arr[211] = 8'b00010010;
		color_arr[212] = 8'b00010010;
		color_arr[213] = 8'b00010010;
		color_arr[214] = 8'b00010010;
		color_arr[215] = 8'b00010010;
		color_arr[216] = 8'b00010010;
		color_arr[217] = 8'b00010010;
		color_arr[218] = 8'b00010010;
		color_arr[219] = 8'b00010010;
		color_arr[220] = 8'b00010010;
		color_arr[221] = 8'b00010010;
		color_arr[222] = 8'b00010010;
		color_arr[223] = 8'b00010010;
		color_arr[224] = 8'b00010010;
		color_arr[225] = 8'b00010010;
		color_arr[226] = 8'b00010010;
		color_arr[227] = 8'b00010010;
		color_arr[228] = 8'b00010010;
		color_arr[229] = 8'b00010010;
		color_arr[230] = 8'b00010010;
		color_arr[231] = 8'b00010010;
		color_arr[232] = 8'b00010010;
		color_arr[233] = 8'b00010010;
		color_arr[234] = 8'b00010010;
		color_arr[235] = 8'b00010010;
		color_arr[236] = 8'b00010010;
		color_arr[237] = 8'b00010010;
		color_arr[238] = 8'b00010010;
		color_arr[239] = 8'b00010010;
		color_arr[240] = 8'b00010010;
		color_arr[241] = 8'b00010010;
		color_arr[242] = 8'b00010010;
		color_arr[243] = 8'b00010010;
		color_arr[244] = 8'b00010010;
		color_arr[245] = 8'b00010010;
		color_arr[246] = 8'b00000000;
		color_arr[247] = 8'b00000000;
		color_arr[248] = 8'b00000000;
		color_arr[249] = 8'b00000000;
		color_arr[250] = 8'b00000000;
		color_arr[251] = 8'b00000000;
		color_arr[252] = 8'b00010010;
		color_arr[253] = 8'b00010010;
		color_arr[254] = 8'b00010010;
		color_arr[255] = 8'b00010010;
		color_arr[256] = 8'b00010010;
		color_arr[257] = 8'b00010010;
		color_arr[258] = 8'b00010010;
		color_arr[259] = 8'b00010010;
		color_arr[260] = 8'b00010010;
		color_arr[261] = 8'b00010010;
		color_arr[262] = 8'b00010010;
		color_arr[263] = 8'b00010010;
		color_arr[264] = 8'b00010010;
		color_arr[265] = 8'b00010010;
		color_arr[266] = 8'b00010010;
		color_arr[267] = 8'b00010010;
		color_arr[268] = 8'b00010010;
		color_arr[269] = 8'b00010010;
		color_arr[270] = 8'b00010010;
		color_arr[271] = 8'b00010010;
		color_arr[272] = 8'b00010010;
		color_arr[273] = 8'b00010010;
		color_arr[274] = 8'b00010010;
		color_arr[275] = 8'b00010010;
		color_arr[276] = 8'b00010010;
		color_arr[277] = 8'b00010010;
		color_arr[278] = 8'b00010010;
		color_arr[279] = 8'b00010010;
		color_arr[280] = 8'b00010010;
		color_arr[281] = 8'b00010010;
		color_arr[282] = 8'b00010010;
		color_arr[283] = 8'b00010010;
		color_arr[284] = 8'b00010010;
		color_arr[285] = 8'b00010010;
		color_arr[286] = 8'b00010010;
		color_arr[287] = 8'b00010010;
		color_arr[288] = 8'b00010010;
		color_arr[289] = 8'b00010010;
		color_arr[290] = 8'b00010010;
		color_arr[291] = 8'b00010010;
		color_arr[292] = 8'b00010010;
		color_arr[293] = 8'b00010010;
		color_arr[294] = 8'b00010010;
		color_arr[295] = 8'b00010010;
		color_arr[296] = 8'b00010010;
		color_arr[297] = 8'b00010010;
		color_arr[298] = 8'b00010010;
		color_arr[299] = 8'b00010010;
		color_arr[300] = 8'b00010010;
		color_arr[301] = 8'b00010010;
		color_arr[302] = 8'b00010010;
		color_arr[303] = 8'b00010010;
		color_arr[304] = 8'b00010010;
		color_arr[305] = 8'b00010010;
		color_arr[306] = 8'b00010010;
		color_arr[307] = 8'b00010010;
		color_arr[308] = 8'b00000000;
		color_arr[309] = 8'b00000000;
		color_arr[310] = 8'b00000000;
		color_arr[311] = 8'b00000000;
		color_arr[312] = 8'b00000000;
		color_arr[313] = 8'b00010010;
		color_arr[314] = 8'b00010010;
		color_arr[315] = 8'b00010010;
		color_arr[316] = 8'b00010010;
		color_arr[317] = 8'b00010010;
		color_arr[318] = 8'b00010010;
		color_arr[319] = 8'b00010010;
		color_arr[320] = 8'b00010010;
		color_arr[321] = 8'b00010010;
		color_arr[322] = 8'b00010010;
		color_arr[323] = 8'b00010010;
		color_arr[324] = 8'b00010010;
		color_arr[325] = 8'b00010010;
		color_arr[326] = 8'b00010010;
		color_arr[327] = 8'b00010010;
		color_arr[328] = 8'b00010010;
		color_arr[329] = 8'b00010010;
		color_arr[330] = 8'b00010010;
		color_arr[331] = 8'b00010010;
		color_arr[332] = 8'b00010010;
		color_arr[333] = 8'b00010010;
		color_arr[334] = 8'b00010010;
		color_arr[335] = 8'b00010010;
		color_arr[336] = 8'b00010010;
		color_arr[337] = 8'b00010010;
		color_arr[338] = 8'b00010010;
		color_arr[339] = 8'b00010010;
		color_arr[340] = 8'b00010010;
		color_arr[341] = 8'b00010010;
		color_arr[342] = 8'b00010010;
		color_arr[343] = 8'b00010010;
		color_arr[344] = 8'b00010010;
		color_arr[345] = 8'b00010010;
		color_arr[346] = 8'b00010010;
		color_arr[347] = 8'b00010010;
		color_arr[348] = 8'b00010010;
		color_arr[349] = 8'b00010010;
		color_arr[350] = 8'b00010010;
		color_arr[351] = 8'b00010010;
		color_arr[352] = 8'b00010010;
		color_arr[353] = 8'b00010010;
		color_arr[354] = 8'b00010010;
		color_arr[355] = 8'b00010010;
		color_arr[356] = 8'b00010010;
		color_arr[357] = 8'b00010010;
		color_arr[358] = 8'b00010010;
		color_arr[359] = 8'b00010010;
		color_arr[360] = 8'b00010010;
		color_arr[361] = 8'b00010010;
		color_arr[362] = 8'b00010010;
		color_arr[363] = 8'b00010010;
		color_arr[364] = 8'b00010010;
		color_arr[365] = 8'b00010010;
		color_arr[366] = 8'b00010010;
		color_arr[367] = 8'b00010010;
		color_arr[368] = 8'b00010010;
		color_arr[369] = 8'b00010010;
		color_arr[370] = 8'b00000000;
		color_arr[371] = 8'b00000000;
		color_arr[372] = 8'b00000000;
		color_arr[373] = 8'b00000000;
		color_arr[374] = 8'b00000000;
		color_arr[375] = 8'b00010010;
		color_arr[376] = 8'b00010010;
		color_arr[377] = 8'b00010010;
		color_arr[378] = 8'b00010010;
		color_arr[379] = 8'b00010010;
		color_arr[380] = 8'b00010010;
		color_arr[381] = 8'b00010010;
		color_arr[382] = 8'b00010010;
		color_arr[383] = 8'b00010010;
		color_arr[384] = 8'b00010010;
		color_arr[385] = 8'b00010010;
		color_arr[386] = 8'b00010010;
		color_arr[387] = 8'b00010010;
		color_arr[388] = 8'b00010010;
		color_arr[389] = 8'b00010010;
		color_arr[390] = 8'b00010010;
		color_arr[391] = 8'b00010010;
		color_arr[392] = 8'b00010010;
		color_arr[393] = 8'b00010010;
		color_arr[394] = 8'b00010010;
		color_arr[395] = 8'b00010010;
		color_arr[396] = 8'b00010010;
		color_arr[397] = 8'b00010010;
		color_arr[398] = 8'b00010010;
		color_arr[399] = 8'b00010010;
		color_arr[400] = 8'b00010010;
		color_arr[401] = 8'b00010010;
		color_arr[402] = 8'b00010010;
		color_arr[403] = 8'b00010010;
		color_arr[404] = 8'b00010010;
		color_arr[405] = 8'b00010010;
		color_arr[406] = 8'b00010010;
		color_arr[407] = 8'b00010010;
		color_arr[408] = 8'b00010010;
		color_arr[409] = 8'b00010010;
		color_arr[410] = 8'b00010010;
		color_arr[411] = 8'b00010010;
		color_arr[412] = 8'b00010010;
		color_arr[413] = 8'b00010010;
		color_arr[414] = 8'b00010010;
		color_arr[415] = 8'b00010010;
		color_arr[416] = 8'b00010010;
		color_arr[417] = 8'b00010010;
		color_arr[418] = 8'b00010010;
		color_arr[419] = 8'b00010010;
		color_arr[420] = 8'b00010010;
		color_arr[421] = 8'b00010010;
		color_arr[422] = 8'b00010010;
		color_arr[423] = 8'b00010010;
		color_arr[424] = 8'b00010010;
		color_arr[425] = 8'b00010010;
		color_arr[426] = 8'b00010010;
		color_arr[427] = 8'b00010010;
		color_arr[428] = 8'b00010010;
		color_arr[429] = 8'b00010010;
		color_arr[430] = 8'b00010010;
		color_arr[431] = 8'b00010010;
		color_arr[432] = 8'b00000000;
		color_arr[433] = 8'b00000000;
		color_arr[434] = 8'b00000000;
		color_arr[435] = 8'b00000000;
		color_arr[436] = 8'b00000000;
		color_arr[437] = 8'b00010010;
		color_arr[438] = 8'b00010010;
		color_arr[439] = 8'b00010010;
		color_arr[440] = 8'b00010010;
		color_arr[441] = 8'b00010010;
		color_arr[442] = 8'b00010010;
		color_arr[443] = 8'b00010010;
		color_arr[444] = 8'b00010010;
		color_arr[445] = 8'b00010010;
		color_arr[446] = 8'b00010010;
		color_arr[447] = 8'b00010010;
		color_arr[448] = 8'b00010010;
		color_arr[449] = 8'b00010010;
		color_arr[450] = 8'b00010010;
		color_arr[451] = 8'b00010010;
		color_arr[452] = 8'b00010010;
		color_arr[453] = 8'b00010010;
		color_arr[454] = 8'b00010010;
		color_arr[455] = 8'b00010010;
		color_arr[456] = 8'b00010010;
		color_arr[457] = 8'b00010010;
		color_arr[458] = 8'b00010010;
		color_arr[459] = 8'b00010010;
		color_arr[460] = 8'b00010010;
		color_arr[461] = 8'b00010010;
		color_arr[462] = 8'b00010010;
		color_arr[463] = 8'b00010010;
		color_arr[464] = 8'b00010010;
		color_arr[465] = 8'b00010010;
		color_arr[466] = 8'b00010010;
		color_arr[467] = 8'b00010010;
		color_arr[468] = 8'b00010010;
		color_arr[469] = 8'b00010010;
		color_arr[470] = 8'b00010010;
		color_arr[471] = 8'b00010010;
		color_arr[472] = 8'b00010010;
		color_arr[473] = 8'b00010010;
		color_arr[474] = 8'b00010010;
		color_arr[475] = 8'b00010010;
		color_arr[476] = 8'b00010010;
		color_arr[477] = 8'b00010010;
		color_arr[478] = 8'b00010010;
		color_arr[479] = 8'b00010010;
		color_arr[480] = 8'b00010010;
		color_arr[481] = 8'b00010010;
		color_arr[482] = 8'b00010010;
		color_arr[483] = 8'b00010010;
		color_arr[484] = 8'b00010010;
		color_arr[485] = 8'b00010010;
		color_arr[486] = 8'b00010010;
		color_arr[487] = 8'b00010010;
		color_arr[488] = 8'b00010010;
		color_arr[489] = 8'b00010010;
		color_arr[490] = 8'b00010010;
		color_arr[491] = 8'b00010010;
		color_arr[492] = 8'b00010010;
		color_arr[493] = 8'b00010010;
		color_arr[494] = 8'b00000000;
		color_arr[495] = 8'b00000000;
		color_arr[496] = 8'b00000000;
		color_arr[497] = 8'b00000000;
		color_arr[498] = 8'b00000000;
		color_arr[499] = 8'b00010010;
		color_arr[500] = 8'b00010010;
		color_arr[501] = 8'b00010010;
		color_arr[502] = 8'b00010010;
		color_arr[503] = 8'b00010010;
		color_arr[504] = 8'b00010010;
		color_arr[505] = 8'b00010010;
		color_arr[506] = 8'b00010010;
		color_arr[507] = 8'b00010010;
		color_arr[508] = 8'b00010010;
		color_arr[509] = 8'b00010010;
		color_arr[510] = 8'b00010010;
		color_arr[511] = 8'b00010010;
		color_arr[512] = 8'b00010010;
		color_arr[513] = 8'b00010010;
		color_arr[514] = 8'b00010010;
		color_arr[515] = 8'b00010010;
		color_arr[516] = 8'b00010010;
		color_arr[517] = 8'b00010010;
		color_arr[518] = 8'b00010010;
		color_arr[519] = 8'b00010010;
		color_arr[520] = 8'b00000010;
		color_arr[521] = 8'b00000010;
		color_arr[522] = 8'b00000010;
		color_arr[523] = 8'b00000010;
		color_arr[524] = 8'b00000010;
		color_arr[525] = 8'b00000010;
		color_arr[526] = 8'b00000010;
		color_arr[527] = 8'b00000010;
		color_arr[528] = 8'b00000010;
		color_arr[529] = 8'b00000010;
		color_arr[530] = 8'b00000010;
		color_arr[531] = 8'b00000010;
		color_arr[532] = 8'b00000010;
		color_arr[533] = 8'b00000010;
		color_arr[534] = 8'b00000010;
		color_arr[535] = 8'b00000010;
		color_arr[536] = 8'b00000010;
		color_arr[537] = 8'b00000010;
		color_arr[538] = 8'b00000010;
		color_arr[539] = 8'b00000010;
		color_arr[540] = 8'b00000010;
		color_arr[541] = 8'b00000010;
		color_arr[542] = 8'b00000010;
		color_arr[543] = 8'b00000010;
		color_arr[544] = 8'b00000010;
		color_arr[545] = 8'b00000010;
		color_arr[546] = 8'b00000010;
		color_arr[547] = 8'b00000010;
		color_arr[548] = 8'b00000010;
		color_arr[549] = 8'b00000010;
		color_arr[550] = 8'b00010010;
		color_arr[551] = 8'b00010010;
		color_arr[552] = 8'b00010010;
		color_arr[553] = 8'b00010010;
		color_arr[554] = 8'b00010010;
		color_arr[555] = 8'b00010010;
		color_arr[556] = 8'b00000000;
		color_arr[557] = 8'b00000000;
		color_arr[558] = 8'b00000000;
		color_arr[559] = 8'b00000000;
		color_arr[560] = 8'b00000000;
		color_arr[561] = 8'b00010010;
		color_arr[562] = 8'b00010010;
		color_arr[563] = 8'b00010010;
		color_arr[564] = 8'b00010010;
		color_arr[565] = 8'b00010010;
		color_arr[566] = 8'b00010010;
		color_arr[567] = 8'b00010010;
		color_arr[568] = 8'b00010010;
		color_arr[569] = 8'b00010010;
		color_arr[570] = 8'b00010010;
		color_arr[571] = 8'b00010010;
		color_arr[572] = 8'b00010010;
		color_arr[573] = 8'b00010010;
		color_arr[574] = 8'b00010010;
		color_arr[575] = 8'b00010010;
		color_arr[576] = 8'b00010010;
		color_arr[577] = 8'b00010010;
		color_arr[578] = 8'b00010010;
		color_arr[579] = 8'b00010010;
		color_arr[580] = 8'b00010010;
		color_arr[581] = 8'b00010010;
		color_arr[582] = 8'b00010010;
		color_arr[583] = 8'b00010010;
		color_arr[584] = 8'b00000010;
		color_arr[585] = 8'b00000010;
		color_arr[586] = 8'b00000010;
		color_arr[587] = 8'b00000010;
		color_arr[588] = 8'b00000010;
		color_arr[589] = 8'b00000010;
		color_arr[590] = 8'b00000010;
		color_arr[591] = 8'b00000010;
		color_arr[592] = 8'b00000010;
		color_arr[593] = 8'b00000010;
		color_arr[594] = 8'b00000010;
		color_arr[595] = 8'b00000010;
		color_arr[596] = 8'b00000010;
		color_arr[597] = 8'b00000010;
		color_arr[598] = 8'b00000010;
		color_arr[599] = 8'b00000010;
		color_arr[600] = 8'b00000010;
		color_arr[601] = 8'b00000010;
		color_arr[602] = 8'b00000010;
		color_arr[603] = 8'b00000010;
		color_arr[604] = 8'b00000010;
		color_arr[605] = 8'b00000010;
		color_arr[606] = 8'b00000010;
		color_arr[607] = 8'b00000010;
		color_arr[608] = 8'b00000010;
		color_arr[609] = 8'b00000010;
		color_arr[610] = 8'b00000010;
		color_arr[611] = 8'b00000010;
		color_arr[612] = 8'b00000010;
		color_arr[613] = 8'b00000010;
		color_arr[614] = 8'b00010010;
		color_arr[615] = 8'b00010010;
		color_arr[616] = 8'b00010010;
		color_arr[617] = 8'b00010010;
		color_arr[618] = 8'b00010010;
		color_arr[619] = 8'b00000000;
		color_arr[620] = 8'b00000000;
		color_arr[621] = 8'b00000000;
		color_arr[622] = 8'b00000000;
		color_arr[623] = 8'b00010010;
		color_arr[624] = 8'b00010010;
		color_arr[625] = 8'b00010010;
		color_arr[626] = 8'b00010010;
		color_arr[627] = 8'b00010010;
		color_arr[628] = 8'b00010010;
		color_arr[629] = 8'b00010010;
		color_arr[630] = 8'b00010010;
		color_arr[631] = 8'b00010010;
		color_arr[632] = 8'b00010010;
		color_arr[633] = 8'b00010010;
		color_arr[634] = 8'b00010010;
		color_arr[635] = 8'b00010010;
		color_arr[636] = 8'b00010010;
		color_arr[637] = 8'b00010010;
		color_arr[638] = 8'b00010010;
		color_arr[639] = 8'b00010010;
		color_arr[640] = 8'b00010010;
		color_arr[641] = 8'b00010010;
		color_arr[642] = 8'b00010010;
		color_arr[643] = 8'b00010010;
		color_arr[644] = 8'b00010010;
		color_arr[645] = 8'b00010010;
		color_arr[646] = 8'b00010010;
		color_arr[647] = 8'b00010010;
		color_arr[648] = 8'b00000010;
		color_arr[649] = 8'b00000010;
		color_arr[650] = 8'b00000010;
		color_arr[651] = 8'b00000010;
		color_arr[652] = 8'b00000010;
		color_arr[653] = 8'b00000010;
		color_arr[654] = 8'b00000010;
		color_arr[655] = 8'b00000010;
		color_arr[656] = 8'b00000010;
		color_arr[657] = 8'b00000010;
		color_arr[658] = 8'b00000010;
		color_arr[659] = 8'b00000010;
		color_arr[660] = 8'b00000010;
		color_arr[661] = 8'b00000010;
		color_arr[662] = 8'b00000010;
		color_arr[663] = 8'b00000010;
		color_arr[664] = 8'b00000010;
		color_arr[665] = 8'b00000010;
		color_arr[666] = 8'b00000010;
		color_arr[667] = 8'b00000010;
		color_arr[668] = 8'b00000010;
		color_arr[669] = 8'b00000010;
		color_arr[670] = 8'b00000010;
		color_arr[671] = 8'b00000010;
		color_arr[672] = 8'b00000010;
		color_arr[673] = 8'b00000010;
		color_arr[674] = 8'b00000010;
		color_arr[675] = 8'b00000010;
		color_arr[676] = 8'b00000010;
		color_arr[677] = 8'b00000010;
		color_arr[678] = 8'b00010010;
		color_arr[679] = 8'b00010010;
		color_arr[680] = 8'b00010010;
		color_arr[681] = 8'b00000000;
		color_arr[682] = 8'b00000000;
		color_arr[683] = 8'b00000000;
		color_arr[684] = 8'b00000000;
		color_arr[685] = 8'b00010010;
		color_arr[686] = 8'b00010010;
		color_arr[687] = 8'b00010010;
		color_arr[688] = 8'b00010010;
		color_arr[689] = 8'b00010010;
		color_arr[690] = 8'b00010010;
		color_arr[691] = 8'b00010010;
		color_arr[692] = 8'b00010010;
		color_arr[693] = 8'b00010010;
		color_arr[694] = 8'b00010010;
		color_arr[695] = 8'b00010010;
		color_arr[696] = 8'b00010010;
		color_arr[697] = 8'b00010010;
		color_arr[698] = 8'b00010010;
		color_arr[699] = 8'b00010010;
		color_arr[700] = 8'b00010010;
		color_arr[701] = 8'b00010010;
		color_arr[702] = 8'b00010010;
		color_arr[703] = 8'b00010010;
		color_arr[704] = 8'b00010010;
		color_arr[705] = 8'b00010010;
		color_arr[706] = 8'b00010010;
		color_arr[707] = 8'b00010010;
		color_arr[708] = 8'b00010010;
		color_arr[709] = 8'b00010010;
		color_arr[710] = 8'b00010010;
		color_arr[711] = 8'b00010010;
		color_arr[712] = 8'b00000010;
		color_arr[713] = 8'b00000010;
		color_arr[714] = 8'b00000010;
		color_arr[715] = 8'b00000010;
		color_arr[716] = 8'b00000010;
		color_arr[717] = 8'b00000010;
		color_arr[718] = 8'b00000010;
		color_arr[719] = 8'b00000010;
		color_arr[720] = 8'b00000010;
		color_arr[721] = 8'b00000010;
		color_arr[722] = 8'b00000010;
		color_arr[723] = 8'b00000010;
		color_arr[724] = 8'b00000010;
		color_arr[725] = 8'b00000010;
		color_arr[726] = 8'b00000010;
		color_arr[727] = 8'b00000010;
		color_arr[728] = 8'b00000010;
		color_arr[729] = 8'b00000010;
		color_arr[730] = 8'b00000010;
		color_arr[731] = 8'b00000010;
		color_arr[732] = 8'b00000010;
		color_arr[733] = 8'b00000010;
		color_arr[734] = 8'b00000010;
		color_arr[735] = 8'b00000010;
		color_arr[736] = 8'b00000010;
		color_arr[737] = 8'b00000010;
		color_arr[738] = 8'b00000010;
		color_arr[739] = 8'b00000010;
		color_arr[740] = 8'b00000010;
		color_arr[741] = 8'b00000010;
		color_arr[742] = 8'b00010010;
		color_arr[743] = 8'b00010010;
		color_arr[744] = 8'b00000000;
		color_arr[745] = 8'b00000000;
		color_arr[746] = 8'b00000000;
		color_arr[747] = 8'b00000000;
		color_arr[748] = 8'b00010010;
		color_arr[749] = 8'b00010010;
		color_arr[750] = 8'b00010010;
		color_arr[751] = 8'b00010010;
		color_arr[752] = 8'b00010010;
		color_arr[753] = 8'b00010010;
		color_arr[754] = 8'b00010010;
		color_arr[755] = 8'b00010010;
		color_arr[756] = 8'b00010010;
		color_arr[757] = 8'b00010010;
		color_arr[758] = 8'b00010010;
		color_arr[759] = 8'b00010010;
		color_arr[760] = 8'b00010010;
		color_arr[761] = 8'b00010010;
		color_arr[762] = 8'b00010010;
		color_arr[763] = 8'b00010010;
		color_arr[764] = 8'b00010010;
		color_arr[765] = 8'b00010010;
		color_arr[766] = 8'b00010010;
		color_arr[767] = 8'b00010010;
		color_arr[768] = 8'b00010010;
		color_arr[769] = 8'b00010010;
		color_arr[770] = 8'b00010010;
		color_arr[771] = 8'b00010010;
		color_arr[772] = 8'b00010010;
		color_arr[773] = 8'b00010010;
		color_arr[774] = 8'b00010010;
		color_arr[775] = 8'b00010010;
		color_arr[776] = 8'b00000010;
		color_arr[777] = 8'b00000010;
		color_arr[778] = 8'b00000010;
		color_arr[779] = 8'b00000010;
		color_arr[780] = 8'b00000010;
		color_arr[781] = 8'b00000010;
		color_arr[782] = 8'b00000010;
		color_arr[783] = 8'b00000010;
		color_arr[784] = 8'b00000010;
		color_arr[785] = 8'b00000010;
		color_arr[786] = 8'b00000010;
		color_arr[787] = 8'b00000010;
		color_arr[788] = 8'b00000010;
		color_arr[789] = 8'b00000010;
		color_arr[790] = 8'b00000010;
		color_arr[791] = 8'b00000010;
		color_arr[792] = 8'b00000010;
		color_arr[793] = 8'b00000010;
		color_arr[794] = 8'b00000010;
		color_arr[795] = 8'b00000010;
		color_arr[796] = 8'b00000010;
		color_arr[797] = 8'b00000010;
		color_arr[798] = 8'b00000010;
		color_arr[799] = 8'b00000010;
		color_arr[800] = 8'b00000010;
		color_arr[801] = 8'b00000010;
		color_arr[802] = 8'b00000010;
		color_arr[803] = 8'b00000010;
		color_arr[804] = 8'b00000010;
		color_arr[805] = 8'b00000010;
		color_arr[806] = 8'b00010010;
		color_arr[807] = 8'b00000000;
		color_arr[808] = 8'b00000000;
		color_arr[809] = 8'b00000000;
		color_arr[810] = 8'b00010010;
		color_arr[811] = 8'b00010010;
		color_arr[812] = 8'b00010010;
		color_arr[813] = 8'b00010010;
		color_arr[814] = 8'b00010010;
		color_arr[815] = 8'b00010010;
		color_arr[816] = 8'b00010010;
		color_arr[817] = 8'b00010010;
		color_arr[818] = 8'b00010010;
		color_arr[819] = 8'b00010010;
		color_arr[820] = 8'b00010010;
		color_arr[821] = 8'b00010010;
		color_arr[822] = 8'b00010010;
		color_arr[823] = 8'b00010010;
		color_arr[824] = 8'b00010010;
		color_arr[825] = 8'b00010010;
		color_arr[826] = 8'b00010010;
		color_arr[827] = 8'b00010010;
		color_arr[828] = 8'b00010010;
		color_arr[829] = 8'b00010010;
		color_arr[830] = 8'b00010010;
		color_arr[831] = 8'b00010010;
		color_arr[832] = 8'b00010010;
		color_arr[833] = 8'b00010010;
		color_arr[834] = 8'b00010010;
		color_arr[835] = 8'b00010010;
		color_arr[836] = 8'b00010010;
		color_arr[837] = 8'b00010010;
		color_arr[838] = 8'b00010010;
		color_arr[839] = 8'b00010010;
		color_arr[840] = 8'b00000010;
		color_arr[841] = 8'b00000010;
		color_arr[842] = 8'b00000010;
		color_arr[843] = 8'b00000010;
		color_arr[844] = 8'b00000010;
		color_arr[845] = 8'b00000010;
		color_arr[846] = 8'b00000010;
		color_arr[847] = 8'b00000010;
		color_arr[848] = 8'b00000010;
		color_arr[849] = 8'b00000010;
		color_arr[850] = 8'b00000010;
		color_arr[851] = 8'b00000010;
		color_arr[852] = 8'b00000010;
		color_arr[853] = 8'b00000010;
		color_arr[854] = 8'b00000010;
		color_arr[855] = 8'b00000010;
		color_arr[856] = 8'b00000010;
		color_arr[857] = 8'b00000010;
		color_arr[858] = 8'b00000010;
		color_arr[859] = 8'b00000010;
		color_arr[860] = 8'b00000010;
		color_arr[861] = 8'b00000010;
		color_arr[862] = 8'b00000010;
		color_arr[863] = 8'b00000010;
		color_arr[864] = 8'b00000010;
		color_arr[865] = 8'b00000010;
		color_arr[866] = 8'b00000010;
		color_arr[867] = 8'b00000010;
		color_arr[868] = 8'b00000010;
		color_arr[869] = 8'b00000010;
		color_arr[870] = 8'b00000000;
		color_arr[871] = 8'b00000000;
		color_arr[872] = 8'b00000000;
		color_arr[873] = 8'b00010010;
		color_arr[874] = 8'b00010010;
		color_arr[875] = 8'b00010010;
		color_arr[876] = 8'b00010010;
		color_arr[877] = 8'b00010010;
		color_arr[878] = 8'b00010010;
		color_arr[879] = 8'b00010010;
		color_arr[880] = 8'b00010010;
		color_arr[881] = 8'b00010010;
		color_arr[882] = 8'b00010010;
		color_arr[883] = 8'b00010010;
		color_arr[884] = 8'b00010010;
		color_arr[885] = 8'b00010010;
		color_arr[886] = 8'b00010010;
		color_arr[887] = 8'b00010010;
		color_arr[888] = 8'b00010010;
		color_arr[889] = 8'b00010010;
		color_arr[890] = 8'b00010010;
		color_arr[891] = 8'b00010010;
		color_arr[892] = 8'b00010010;
		color_arr[893] = 8'b00010010;
		color_arr[894] = 8'b00010010;
		color_arr[895] = 8'b00010010;
		color_arr[896] = 8'b00010010;
		color_arr[897] = 8'b00010010;
		color_arr[898] = 8'b00010010;
		color_arr[899] = 8'b00010010;
		color_arr[900] = 8'b00010010;
		color_arr[901] = 8'b00010010;
		color_arr[902] = 8'b00010010;
		color_arr[903] = 8'b00010010;
		color_arr[904] = 8'b00000010;
		color_arr[905] = 8'b00000010;
		color_arr[906] = 8'b00000010;
		color_arr[907] = 8'b00000010;
		color_arr[908] = 8'b00000010;
		color_arr[909] = 8'b00000010;
		color_arr[910] = 8'b00000010;
		color_arr[911] = 8'b00000010;
		color_arr[912] = 8'b00000010;
		color_arr[913] = 8'b00000010;
		color_arr[914] = 8'b00000010;
		color_arr[915] = 8'b00000010;
		color_arr[916] = 8'b00000010;
		color_arr[917] = 8'b00000010;
		color_arr[918] = 8'b00000010;
		color_arr[919] = 8'b00000010;
		color_arr[920] = 8'b00000010;
		color_arr[921] = 8'b00000010;
		color_arr[922] = 8'b00000010;
		color_arr[923] = 8'b00000010;
		color_arr[924] = 8'b00000010;
		color_arr[925] = 8'b00000010;
		color_arr[926] = 8'b00000010;
		color_arr[927] = 8'b00000010;
		color_arr[928] = 8'b00000010;
		color_arr[929] = 8'b00000010;
		color_arr[930] = 8'b00000010;
		color_arr[931] = 8'b00000010;
		color_arr[932] = 8'b00000000;
		color_arr[933] = 8'b00000000;
		color_arr[934] = 8'b00000000;
		color_arr[935] = 8'b00000000;
		color_arr[936] = 8'b00010010;
		color_arr[937] = 8'b00010010;
		color_arr[938] = 8'b00010010;
		color_arr[939] = 8'b00010010;
		color_arr[940] = 8'b00010010;
		color_arr[941] = 8'b00010010;
		color_arr[942] = 8'b00010010;
		color_arr[943] = 8'b00010010;
		color_arr[944] = 8'b00010010;
		color_arr[945] = 8'b00010010;
		color_arr[946] = 8'b00010010;
		color_arr[947] = 8'b00010010;
		color_arr[948] = 8'b00010010;
		color_arr[949] = 8'b00010010;
		color_arr[950] = 8'b00010010;
		color_arr[951] = 8'b00010010;
		color_arr[952] = 8'b00010010;
		color_arr[953] = 8'b00010010;
		color_arr[954] = 8'b00010010;
		color_arr[955] = 8'b00010010;
		color_arr[956] = 8'b00010010;
		color_arr[957] = 8'b00010010;
		color_arr[958] = 8'b00010010;
		color_arr[959] = 8'b00010010;
		color_arr[960] = 8'b00010010;
		color_arr[961] = 8'b00010010;
		color_arr[962] = 8'b00010010;
		color_arr[963] = 8'b00010010;
		color_arr[964] = 8'b00010010;
		color_arr[965] = 8'b00010010;
		color_arr[966] = 8'b00010010;
		color_arr[967] = 8'b00010010;
		color_arr[968] = 8'b00000010;
		color_arr[969] = 8'b00000010;
		color_arr[970] = 8'b00000010;
		color_arr[971] = 8'b00000010;
		color_arr[972] = 8'b00000010;
		color_arr[973] = 8'b00000010;
		color_arr[974] = 8'b00000010;
		color_arr[975] = 8'b00000010;
		color_arr[976] = 8'b00000010;
		color_arr[977] = 8'b00000010;
		color_arr[978] = 8'b00000010;
		color_arr[979] = 8'b00000010;
		color_arr[980] = 8'b00000010;
		color_arr[981] = 8'b00000010;
		color_arr[982] = 8'b00000010;
		color_arr[983] = 8'b00000010;
		color_arr[984] = 8'b00000010;
		color_arr[985] = 8'b00000010;
		color_arr[986] = 8'b00000010;
		color_arr[987] = 8'b00000010;
		color_arr[988] = 8'b00000010;
		color_arr[989] = 8'b00000010;
		color_arr[990] = 8'b00000010;
		color_arr[991] = 8'b00000010;
		color_arr[992] = 8'b00000010;
		color_arr[993] = 8'b00000010;
		color_arr[994] = 8'b00000010;
		color_arr[995] = 8'b00000000;
		color_arr[996] = 8'b00000000;
		color_arr[997] = 8'b00000000;
		color_arr[998] = 8'b00000000;
		color_arr[999] = 8'b00010010;
		color_arr[1000] = 8'b00010010;
		color_arr[1001] = 8'b00010010;
		color_arr[1002] = 8'b00010010;
		color_arr[1003] = 8'b00010010;
		color_arr[1004] = 8'b00010010;
		color_arr[1005] = 8'b00010010;
		color_arr[1006] = 8'b00010010;
		color_arr[1007] = 8'b00010010;
		color_arr[1008] = 8'b00010010;
		color_arr[1009] = 8'b00010010;
		color_arr[1010] = 8'b00010010;
		color_arr[1011] = 8'b00010010;
		color_arr[1012] = 8'b00010010;
		color_arr[1013] = 8'b00010010;
		color_arr[1014] = 8'b00010010;
		color_arr[1015] = 8'b00010010;
		color_arr[1016] = 8'b00010010;
		color_arr[1017] = 8'b00010010;
		color_arr[1018] = 8'b00010010;
		color_arr[1019] = 8'b00010010;
		color_arr[1020] = 8'b00010010;
		color_arr[1021] = 8'b00010010;
		color_arr[1022] = 8'b00010010;
		color_arr[1023] = 8'b00010010;
		color_arr[1024] = 8'b00010010;
		color_arr[1025] = 8'b00010010;
		color_arr[1026] = 8'b00010010;
		color_arr[1027] = 8'b00010010;
		color_arr[1028] = 8'b00010010;
		color_arr[1029] = 8'b00010010;
		color_arr[1030] = 8'b00010010;
		color_arr[1031] = 8'b00010010;
		color_arr[1032] = 8'b00000010;
		color_arr[1033] = 8'b00000010;
		color_arr[1034] = 8'b00000010;
		color_arr[1035] = 8'b00000010;
		color_arr[1036] = 8'b00000010;
		color_arr[1037] = 8'b00000010;
		color_arr[1038] = 8'b00000010;
		color_arr[1039] = 8'b00000010;
		color_arr[1040] = 8'b00000010;
		color_arr[1041] = 8'b00000010;
		color_arr[1042] = 8'b00000010;
		color_arr[1043] = 8'b00000010;
		color_arr[1044] = 8'b00000010;
		color_arr[1045] = 8'b00000010;
		color_arr[1046] = 8'b00000010;
		color_arr[1047] = 8'b00000010;
		color_arr[1048] = 8'b00000010;
		color_arr[1049] = 8'b00000010;
		color_arr[1050] = 8'b00000010;
		color_arr[1051] = 8'b00000010;
		color_arr[1052] = 8'b00000010;
		color_arr[1053] = 8'b00000010;
		color_arr[1054] = 8'b00000010;
		color_arr[1055] = 8'b00000010;
		color_arr[1056] = 8'b00000010;
		color_arr[1057] = 8'b00000010;
		color_arr[1058] = 8'b00000000;
		color_arr[1059] = 8'b00000000;
		color_arr[1060] = 8'b00000000;
		color_arr[1061] = 8'b00000010;
		color_arr[1062] = 8'b00010010;
		color_arr[1063] = 8'b00010010;
		color_arr[1064] = 8'b00010010;
		color_arr[1065] = 8'b00010010;
		color_arr[1066] = 8'b00010010;
		color_arr[1067] = 8'b00010010;
		color_arr[1068] = 8'b00010010;
		color_arr[1069] = 8'b00010010;
		color_arr[1070] = 8'b00010010;
		color_arr[1071] = 8'b00010010;
		color_arr[1072] = 8'b00010010;
		color_arr[1073] = 8'b00010010;
		color_arr[1074] = 8'b00010010;
		color_arr[1075] = 8'b00010010;
		color_arr[1076] = 8'b00010010;
		color_arr[1077] = 8'b00010010;
		color_arr[1078] = 8'b00010010;
		color_arr[1079] = 8'b00010010;
		color_arr[1080] = 8'b00010010;
		color_arr[1081] = 8'b00010010;
		color_arr[1082] = 8'b00010010;
		color_arr[1083] = 8'b00010010;
		color_arr[1084] = 8'b00010010;
		color_arr[1085] = 8'b00010010;
		color_arr[1086] = 8'b00010010;
		color_arr[1087] = 8'b00010010;
		color_arr[1088] = 8'b00010010;
		color_arr[1089] = 8'b00010010;
		color_arr[1090] = 8'b00010010;
		color_arr[1091] = 8'b00010010;
		color_arr[1092] = 8'b00010010;
		color_arr[1093] = 8'b00010010;
		color_arr[1094] = 8'b00010010;
		color_arr[1095] = 8'b00010010;
		color_arr[1096] = 8'b00000010;
		color_arr[1097] = 8'b00000010;
		color_arr[1098] = 8'b00000010;
		color_arr[1099] = 8'b00000010;
		color_arr[1100] = 8'b00000010;
		color_arr[1101] = 8'b00000010;
		color_arr[1102] = 8'b00000010;
		color_arr[1103] = 8'b00000010;
		color_arr[1104] = 8'b00000010;
		color_arr[1105] = 8'b00000010;
		color_arr[1106] = 8'b00000010;
		color_arr[1107] = 8'b00000010;
		color_arr[1108] = 8'b00000010;
		color_arr[1109] = 8'b00000010;
		color_arr[1110] = 8'b00000010;
		color_arr[1111] = 8'b00000010;
		color_arr[1112] = 8'b00000010;
		color_arr[1113] = 8'b00000010;
		color_arr[1114] = 8'b00000010;
		color_arr[1115] = 8'b00000010;
		color_arr[1116] = 8'b00000010;
		color_arr[1117] = 8'b00000010;
		color_arr[1118] = 8'b00000010;
		color_arr[1119] = 8'b00000010;
		color_arr[1120] = 8'b00000010;
		color_arr[1121] = 8'b00000000;
		color_arr[1122] = 8'b00000000;
		color_arr[1123] = 8'b00000000;
		color_arr[1124] = 8'b00000010;
		color_arr[1125] = 8'b00000010;
		color_arr[1126] = 8'b00010010;
		color_arr[1127] = 8'b00010010;
		color_arr[1128] = 8'b00010010;
		color_arr[1129] = 8'b00010010;
		color_arr[1130] = 8'b00010010;
		color_arr[1131] = 8'b00010010;
		color_arr[1132] = 8'b00010010;
		color_arr[1133] = 8'b00010010;
		color_arr[1134] = 8'b00010010;
		color_arr[1135] = 8'b00010010;
		color_arr[1136] = 8'b00010010;
		color_arr[1137] = 8'b00010010;
		color_arr[1138] = 8'b00010010;
		color_arr[1139] = 8'b00010010;
		color_arr[1140] = 8'b00010010;
		color_arr[1141] = 8'b00010010;
		color_arr[1142] = 8'b00010010;
		color_arr[1143] = 8'b00010010;
		color_arr[1144] = 8'b00010010;
		color_arr[1145] = 8'b00010010;
		color_arr[1146] = 8'b00010010;
		color_arr[1147] = 8'b00010010;
		color_arr[1148] = 8'b00010010;
		color_arr[1149] = 8'b00010010;
		color_arr[1150] = 8'b00010010;
		color_arr[1151] = 8'b00010010;
		color_arr[1152] = 8'b00010010;
		color_arr[1153] = 8'b00010010;
		color_arr[1154] = 8'b00010010;
		color_arr[1155] = 8'b00010010;
		color_arr[1156] = 8'b00010010;
		color_arr[1157] = 8'b00010010;
		color_arr[1158] = 8'b00010010;
		color_arr[1159] = 8'b00010010;
		color_arr[1160] = 8'b00000010;
		color_arr[1161] = 8'b00000010;
		color_arr[1162] = 8'b00000010;
		color_arr[1163] = 8'b00000010;
		color_arr[1164] = 8'b00000010;
		color_arr[1165] = 8'b00000010;
		color_arr[1166] = 8'b00000010;
		color_arr[1167] = 8'b00000010;
		color_arr[1168] = 8'b00000010;
		color_arr[1169] = 8'b00000010;
		color_arr[1170] = 8'b00000010;
		color_arr[1171] = 8'b00000010;
		color_arr[1172] = 8'b00000010;
		color_arr[1173] = 8'b00000010;
		color_arr[1174] = 8'b00000010;
		color_arr[1175] = 8'b00000010;
		color_arr[1176] = 8'b00000010;
		color_arr[1177] = 8'b00000010;
		color_arr[1178] = 8'b00000010;
		color_arr[1179] = 8'b00000010;
		color_arr[1180] = 8'b00000010;
		color_arr[1181] = 8'b00000010;
		color_arr[1182] = 8'b00000010;
		color_arr[1183] = 8'b00000010;
		color_arr[1184] = 8'b00000000;
		color_arr[1185] = 8'b00000000;
		color_arr[1186] = 8'b00000000;
		color_arr[1187] = 8'b00000010;
		color_arr[1188] = 8'b00000010;
		color_arr[1189] = 8'b00000010;
		color_arr[1190] = 8'b00010010;
		color_arr[1191] = 8'b00010010;
		color_arr[1192] = 8'b00010010;
		color_arr[1193] = 8'b00010010;
		color_arr[1194] = 8'b00010010;
		color_arr[1195] = 8'b00010010;
		color_arr[1196] = 8'b00010010;
		color_arr[1197] = 8'b00010010;
		color_arr[1198] = 8'b00010010;
		color_arr[1199] = 8'b00010010;
		color_arr[1200] = 8'b00010010;
		color_arr[1201] = 8'b00010010;
		color_arr[1202] = 8'b00010010;
		color_arr[1203] = 8'b00010010;
		color_arr[1204] = 8'b00010010;
		color_arr[1205] = 8'b00010010;
		color_arr[1206] = 8'b00010010;
		color_arr[1207] = 8'b00010010;
		color_arr[1208] = 8'b00010010;
		color_arr[1209] = 8'b00010010;
		color_arr[1210] = 8'b00010010;
		color_arr[1211] = 8'b00010010;
		color_arr[1212] = 8'b00010010;
		color_arr[1213] = 8'b00010010;
		color_arr[1214] = 8'b00010010;
		color_arr[1215] = 8'b00010010;
		color_arr[1216] = 8'b00010010;
		color_arr[1217] = 8'b00010010;
		color_arr[1218] = 8'b00010010;
		color_arr[1219] = 8'b00010010;
		color_arr[1220] = 8'b00010010;
		color_arr[1221] = 8'b00010010;
		color_arr[1222] = 8'b00010010;
		color_arr[1223] = 8'b00010010;
		color_arr[1224] = 8'b00000010;
		color_arr[1225] = 8'b00000010;
		color_arr[1226] = 8'b00000010;
		color_arr[1227] = 8'b00000010;
		color_arr[1228] = 8'b00000010;
		color_arr[1229] = 8'b00000010;
		color_arr[1230] = 8'b00000010;
		color_arr[1231] = 8'b00000010;
		color_arr[1232] = 8'b00000010;
		color_arr[1233] = 8'b00000010;
		color_arr[1234] = 8'b00000010;
		color_arr[1235] = 8'b00000010;
		color_arr[1236] = 8'b00000010;
		color_arr[1237] = 8'b00000010;
		color_arr[1238] = 8'b00000010;
		color_arr[1239] = 8'b00000010;
		color_arr[1240] = 8'b00000010;
		color_arr[1241] = 8'b00000010;
		color_arr[1242] = 8'b00000010;
		color_arr[1243] = 8'b00000010;
		color_arr[1244] = 8'b00000010;
		color_arr[1245] = 8'b00000010;
		color_arr[1246] = 8'b00000010;
		color_arr[1247] = 8'b00000000;
		color_arr[1248] = 8'b00000000;
		color_arr[1249] = 8'b00000000;
		color_arr[1250] = 8'b00000010;
		color_arr[1251] = 8'b00000010;
		color_arr[1252] = 8'b00000010;
		color_arr[1253] = 8'b00000010;
		color_arr[1254] = 8'b00010010;
		color_arr[1255] = 8'b00010010;
		color_arr[1256] = 8'b00010010;
		color_arr[1257] = 8'b00010010;
		color_arr[1258] = 8'b00010010;
		color_arr[1259] = 8'b00010010;
		color_arr[1260] = 8'b00010010;
		color_arr[1261] = 8'b00010010;
		color_arr[1262] = 8'b00010010;
		color_arr[1263] = 8'b00010010;
		color_arr[1264] = 8'b00010010;
		color_arr[1265] = 8'b00010010;
		color_arr[1266] = 8'b00010010;
		color_arr[1267] = 8'b00010010;
		color_arr[1268] = 8'b00010010;
		color_arr[1269] = 8'b00010010;
		color_arr[1270] = 8'b00010010;
		color_arr[1271] = 8'b00010010;
		color_arr[1272] = 8'b00010010;
		color_arr[1273] = 8'b00010010;
		color_arr[1274] = 8'b00010010;
		color_arr[1275] = 8'b00010010;
		color_arr[1276] = 8'b00010010;
		color_arr[1277] = 8'b00010010;
		color_arr[1278] = 8'b00010010;
		color_arr[1279] = 8'b00010010;
		color_arr[1280] = 8'b00010010;
		color_arr[1281] = 8'b00010010;
		color_arr[1282] = 8'b00010010;
		color_arr[1283] = 8'b00010010;
		color_arr[1284] = 8'b00010010;
		color_arr[1285] = 8'b00010010;
		color_arr[1286] = 8'b00010010;
		color_arr[1287] = 8'b00010010;
		color_arr[1288] = 8'b00000010;
		color_arr[1289] = 8'b00000010;
		color_arr[1290] = 8'b00000010;
		color_arr[1291] = 8'b00000010;
		color_arr[1292] = 8'b00000010;
		color_arr[1293] = 8'b00000010;
		color_arr[1294] = 8'b00000010;
		color_arr[1295] = 8'b00000010;
		color_arr[1296] = 8'b00000010;
		color_arr[1297] = 8'b00000010;
		color_arr[1298] = 8'b00000010;
		color_arr[1299] = 8'b00000010;
		color_arr[1300] = 8'b00000010;
		color_arr[1301] = 8'b00000010;
		color_arr[1302] = 8'b00000010;
		color_arr[1303] = 8'b00000010;
		color_arr[1304] = 8'b00000010;
		color_arr[1305] = 8'b00000010;
		color_arr[1306] = 8'b00000010;
		color_arr[1307] = 8'b00000010;
		color_arr[1308] = 8'b00000010;
		color_arr[1309] = 8'b00000010;
		color_arr[1310] = 8'b00000000;
		color_arr[1311] = 8'b00000000;
		color_arr[1312] = 8'b00000000;
		color_arr[1313] = 8'b00000010;
		color_arr[1314] = 8'b00000010;
		color_arr[1315] = 8'b00000010;
		color_arr[1316] = 8'b00000010;
		color_arr[1317] = 8'b00000010;
		color_arr[1318] = 8'b00010010;
		color_arr[1319] = 8'b00010010;
		color_arr[1320] = 8'b00010010;
		color_arr[1321] = 8'b00010010;
		color_arr[1322] = 8'b00010010;
		color_arr[1323] = 8'b00010010;
		color_arr[1324] = 8'b00010010;
		color_arr[1325] = 8'b00010010;
		color_arr[1326] = 8'b00010010;
		color_arr[1327] = 8'b00010010;
		color_arr[1328] = 8'b00010010;
		color_arr[1329] = 8'b00010010;
		color_arr[1330] = 8'b00010010;
		color_arr[1331] = 8'b00010010;
		color_arr[1332] = 8'b00010010;
		color_arr[1333] = 8'b00010010;
		color_arr[1334] = 8'b00010010;
		color_arr[1335] = 8'b00010010;
		color_arr[1336] = 8'b00010010;
		color_arr[1337] = 8'b00010010;
		color_arr[1338] = 8'b00010010;
		color_arr[1339] = 8'b00010010;
		color_arr[1340] = 8'b00010010;
		color_arr[1341] = 8'b00010010;
		color_arr[1342] = 8'b00010010;
		color_arr[1343] = 8'b00010010;
		color_arr[1344] = 8'b00010010;
		color_arr[1345] = 8'b00010010;
		color_arr[1346] = 8'b00010010;
		color_arr[1347] = 8'b00010010;
		color_arr[1348] = 8'b00010010;
		color_arr[1349] = 8'b00010010;
		color_arr[1350] = 8'b00010010;
		color_arr[1351] = 8'b00010010;
		color_arr[1352] = 8'b00000010;
		color_arr[1353] = 8'b00000010;
		color_arr[1354] = 8'b00000010;
		color_arr[1355] = 8'b00000010;
		color_arr[1356] = 8'b00000010;
		color_arr[1357] = 8'b00000010;
		color_arr[1358] = 8'b00000010;
		color_arr[1359] = 8'b00000010;
		color_arr[1360] = 8'b00000010;
		color_arr[1361] = 8'b00000010;
		color_arr[1362] = 8'b00000010;
		color_arr[1363] = 8'b00000010;
		color_arr[1364] = 8'b00000010;
		color_arr[1365] = 8'b00000010;
		color_arr[1366] = 8'b00000010;
		color_arr[1367] = 8'b00000010;
		color_arr[1368] = 8'b00000010;
		color_arr[1369] = 8'b00000010;
		color_arr[1370] = 8'b00000010;
		color_arr[1371] = 8'b00000010;
		color_arr[1372] = 8'b00000010;
		color_arr[1373] = 8'b00000000;
		color_arr[1374] = 8'b00000000;
		color_arr[1375] = 8'b00000000;
		color_arr[1376] = 8'b00000010;
		color_arr[1377] = 8'b00000010;
		color_arr[1378] = 8'b00000010;
		color_arr[1379] = 8'b00000010;
		color_arr[1380] = 8'b00000010;
		color_arr[1381] = 8'b00000010;
		color_arr[1382] = 8'b00010010;
		color_arr[1383] = 8'b00010010;
		color_arr[1384] = 8'b00010010;
		color_arr[1385] = 8'b00010010;
		color_arr[1386] = 8'b00010010;
		color_arr[1387] = 8'b00010010;
		color_arr[1388] = 8'b00010010;
		color_arr[1389] = 8'b00010010;
		color_arr[1390] = 8'b00010010;
		color_arr[1391] = 8'b00010010;
		color_arr[1392] = 8'b00010010;
		color_arr[1393] = 8'b00010010;
		color_arr[1394] = 8'b00010010;
		color_arr[1395] = 8'b00010010;
		color_arr[1396] = 8'b00010010;
		color_arr[1397] = 8'b00010010;
		color_arr[1398] = 8'b00010010;
		color_arr[1399] = 8'b00010010;
		color_arr[1400] = 8'b00010010;
		color_arr[1401] = 8'b00010010;
		color_arr[1402] = 8'b00010010;
		color_arr[1403] = 8'b00010010;
		color_arr[1404] = 8'b00010010;
		color_arr[1405] = 8'b00010010;
		color_arr[1406] = 8'b00010010;
		color_arr[1407] = 8'b00010010;
		color_arr[1408] = 8'b00010010;
		color_arr[1409] = 8'b00010010;
		color_arr[1410] = 8'b00010010;
		color_arr[1411] = 8'b00010010;
		color_arr[1412] = 8'b00010010;
		color_arr[1413] = 8'b00010010;
		color_arr[1414] = 8'b00010010;
		color_arr[1415] = 8'b00010010;
		color_arr[1416] = 8'b00000010;
		color_arr[1417] = 8'b00000010;
		color_arr[1418] = 8'b00000010;
		color_arr[1419] = 8'b00000010;
		color_arr[1420] = 8'b00000010;
		color_arr[1421] = 8'b00000010;
		color_arr[1422] = 8'b00000010;
		color_arr[1423] = 8'b00000010;
		color_arr[1424] = 8'b00000010;
		color_arr[1425] = 8'b00000010;
		color_arr[1426] = 8'b00000010;
		color_arr[1427] = 8'b00000010;
		color_arr[1428] = 8'b00000010;
		color_arr[1429] = 8'b00000010;
		color_arr[1430] = 8'b00000010;
		color_arr[1431] = 8'b00000010;
		color_arr[1432] = 8'b00000010;
		color_arr[1433] = 8'b00000010;
		color_arr[1434] = 8'b00000010;
		color_arr[1435] = 8'b00000010;
		color_arr[1436] = 8'b00000000;
		color_arr[1437] = 8'b00000000;
		color_arr[1438] = 8'b00000000;
		color_arr[1439] = 8'b00000010;
		color_arr[1440] = 8'b00000010;
		color_arr[1441] = 8'b00000010;
		color_arr[1442] = 8'b00000010;
		color_arr[1443] = 8'b00000010;
		color_arr[1444] = 8'b00000010;
		color_arr[1445] = 8'b00000010;
		color_arr[1446] = 8'b00100000;
		color_arr[1447] = 8'b00100000;
		color_arr[1448] = 8'b00100000;
		color_arr[1449] = 8'b00100000;
		color_arr[1450] = 8'b00100000;
		color_arr[1451] = 8'b00100000;
		color_arr[1452] = 8'b00100000;
		color_arr[1453] = 8'b00100000;
		color_arr[1454] = 8'b00100000;
		color_arr[1455] = 8'b00100000;
		color_arr[1456] = 8'b00100000;
		color_arr[1457] = 8'b00100000;
		color_arr[1458] = 8'b00100000;
		color_arr[1459] = 8'b00100000;
		color_arr[1460] = 8'b00100000;
		color_arr[1461] = 8'b00100000;
		color_arr[1462] = 8'b00100000;
		color_arr[1463] = 8'b00100000;
		color_arr[1464] = 8'b00100000;
		color_arr[1465] = 8'b00100000;
		color_arr[1466] = 8'b00100000;
		color_arr[1467] = 8'b00100000;
		color_arr[1468] = 8'b00100000;
		color_arr[1469] = 8'b00100000;
		color_arr[1470] = 8'b00100000;
		color_arr[1471] = 8'b00100000;
		color_arr[1472] = 8'b00010010;
		color_arr[1473] = 8'b00010010;
		color_arr[1474] = 8'b00010010;
		color_arr[1475] = 8'b00010010;
		color_arr[1476] = 8'b00010010;
		color_arr[1477] = 8'b00010010;
		color_arr[1478] = 8'b00010010;
		color_arr[1479] = 8'b00010010;
		color_arr[1480] = 8'b00000010;
		color_arr[1481] = 8'b00000010;
		color_arr[1482] = 8'b00000010;
		color_arr[1483] = 8'b00000010;
		color_arr[1484] = 8'b00000010;
		color_arr[1485] = 8'b00000010;
		color_arr[1486] = 8'b00000010;
		color_arr[1487] = 8'b00000010;
		color_arr[1488] = 8'b00000010;
		color_arr[1489] = 8'b00000010;
		color_arr[1490] = 8'b00000010;
		color_arr[1491] = 8'b00000010;
		color_arr[1492] = 8'b00000010;
		color_arr[1493] = 8'b00000010;
		color_arr[1494] = 8'b00000010;
		color_arr[1495] = 8'b00000010;
		color_arr[1496] = 8'b00000010;
		color_arr[1497] = 8'b00000010;
		color_arr[1498] = 8'b00000010;
		color_arr[1499] = 8'b00000000;
		color_arr[1500] = 8'b00000000;
		color_arr[1501] = 8'b00000000;
		color_arr[1502] = 8'b00000010;
		color_arr[1503] = 8'b00000010;
		color_arr[1504] = 8'b00000010;
		color_arr[1505] = 8'b00000010;
		color_arr[1506] = 8'b00000010;
		color_arr[1507] = 8'b00000010;
		color_arr[1508] = 8'b00000010;
		color_arr[1509] = 8'b00000010;
		color_arr[1510] = 8'b00100000;
		color_arr[1511] = 8'b00100000;
		color_arr[1512] = 8'b00100000;
		color_arr[1513] = 8'b00100000;
		color_arr[1514] = 8'b00100000;
		color_arr[1515] = 8'b00100000;
		color_arr[1516] = 8'b00100000;
		color_arr[1517] = 8'b00100000;
		color_arr[1518] = 8'b00100000;
		color_arr[1519] = 8'b00100000;
		color_arr[1520] = 8'b00100000;
		color_arr[1521] = 8'b00100000;
		color_arr[1522] = 8'b00100000;
		color_arr[1523] = 8'b00100000;
		color_arr[1524] = 8'b00100000;
		color_arr[1525] = 8'b00100000;
		color_arr[1526] = 8'b00100000;
		color_arr[1527] = 8'b00100000;
		color_arr[1528] = 8'b00100000;
		color_arr[1529] = 8'b00100000;
		color_arr[1530] = 8'b00100000;
		color_arr[1531] = 8'b00100000;
		color_arr[1532] = 8'b00100000;
		color_arr[1533] = 8'b00100000;
		color_arr[1534] = 8'b00100000;
		color_arr[1535] = 8'b00100000;
		color_arr[1536] = 8'b00010010;
		color_arr[1537] = 8'b00010010;
		color_arr[1538] = 8'b00010010;
		color_arr[1539] = 8'b00010010;
		color_arr[1540] = 8'b00010010;
		color_arr[1541] = 8'b00010010;
		color_arr[1542] = 8'b00010010;
		color_arr[1543] = 8'b00010010;
		color_arr[1544] = 8'b00000010;
		color_arr[1545] = 8'b00000010;
		color_arr[1546] = 8'b00000010;
		color_arr[1547] = 8'b00000010;
		color_arr[1548] = 8'b00000010;
		color_arr[1549] = 8'b00000010;
		color_arr[1550] = 8'b00000010;
		color_arr[1551] = 8'b00000010;
		color_arr[1552] = 8'b00000010;
		color_arr[1553] = 8'b00000010;
		color_arr[1554] = 8'b00000010;
		color_arr[1555] = 8'b00000010;
		color_arr[1556] = 8'b00000010;
		color_arr[1557] = 8'b00000010;
		color_arr[1558] = 8'b00000010;
		color_arr[1559] = 8'b00000010;
		color_arr[1560] = 8'b00000010;
		color_arr[1561] = 8'b00000010;
		color_arr[1562] = 8'b00000000;
		color_arr[1563] = 8'b00000000;
		color_arr[1564] = 8'b00000000;
		color_arr[1565] = 8'b00000010;
		color_arr[1566] = 8'b00000010;
		color_arr[1567] = 8'b00000010;
		color_arr[1568] = 8'b00000010;
		color_arr[1569] = 8'b00000010;
		color_arr[1570] = 8'b00000010;
		color_arr[1571] = 8'b00000010;
		color_arr[1572] = 8'b00000010;
		color_arr[1573] = 8'b00000010;
		color_arr[1574] = 8'b00100000;
		color_arr[1575] = 8'b00100000;
		color_arr[1576] = 8'b00100000;
		color_arr[1577] = 8'b00100000;
		color_arr[1578] = 8'b00100000;
		color_arr[1579] = 8'b00100000;
		color_arr[1580] = 8'b00100000;
		color_arr[1581] = 8'b00100000;
		color_arr[1582] = 8'b00100000;
		color_arr[1583] = 8'b00100000;
		color_arr[1584] = 8'b00100000;
		color_arr[1585] = 8'b00100000;
		color_arr[1586] = 8'b00100000;
		color_arr[1587] = 8'b00100000;
		color_arr[1588] = 8'b00100000;
		color_arr[1589] = 8'b00100000;
		color_arr[1590] = 8'b00100000;
		color_arr[1591] = 8'b00100000;
		color_arr[1592] = 8'b00100000;
		color_arr[1593] = 8'b00100000;
		color_arr[1594] = 8'b00100000;
		color_arr[1595] = 8'b00100000;
		color_arr[1596] = 8'b00100000;
		color_arr[1597] = 8'b00100000;
		color_arr[1598] = 8'b00100000;
		color_arr[1599] = 8'b00100000;
		color_arr[1600] = 8'b00010010;
		color_arr[1601] = 8'b00010010;
		color_arr[1602] = 8'b00010010;
		color_arr[1603] = 8'b00010010;
		color_arr[1604] = 8'b00010010;
		color_arr[1605] = 8'b00010010;
		color_arr[1606] = 8'b00010010;
		color_arr[1607] = 8'b00010010;
		color_arr[1608] = 8'b00000010;
		color_arr[1609] = 8'b00000010;
		color_arr[1610] = 8'b00000010;
		color_arr[1611] = 8'b00000010;
		color_arr[1612] = 8'b00000010;
		color_arr[1613] = 8'b00000010;
		color_arr[1614] = 8'b00000010;
		color_arr[1615] = 8'b00000010;
		color_arr[1616] = 8'b00000010;
		color_arr[1617] = 8'b00000010;
		color_arr[1618] = 8'b00000010;
		color_arr[1619] = 8'b00000010;
		color_arr[1620] = 8'b00000010;
		color_arr[1621] = 8'b00000010;
		color_arr[1622] = 8'b00000010;
		color_arr[1623] = 8'b00000010;
		color_arr[1624] = 8'b00000010;
		color_arr[1625] = 8'b00000000;
		color_arr[1626] = 8'b00000000;
		color_arr[1627] = 8'b00000000;
		color_arr[1628] = 8'b00000010;
		color_arr[1629] = 8'b00000010;
		color_arr[1630] = 8'b00000010;
		color_arr[1631] = 8'b00000010;
		color_arr[1632] = 8'b00000010;
		color_arr[1633] = 8'b00000010;
		color_arr[1634] = 8'b00000010;
		color_arr[1635] = 8'b00000010;
		color_arr[1636] = 8'b00000010;
		color_arr[1637] = 8'b00000010;
		color_arr[1638] = 8'b00100000;
		color_arr[1639] = 8'b00100000;
		color_arr[1640] = 8'b00100000;
		color_arr[1641] = 8'b00100000;
		color_arr[1642] = 8'b00100000;
		color_arr[1643] = 8'b00100000;
		color_arr[1644] = 8'b00100000;
		color_arr[1645] = 8'b00100000;
		color_arr[1646] = 8'b00100000;
		color_arr[1647] = 8'b00100000;
		color_arr[1648] = 8'b00100000;
		color_arr[1649] = 8'b00100000;
		color_arr[1650] = 8'b00100000;
		color_arr[1651] = 8'b00100000;
		color_arr[1652] = 8'b00100000;
		color_arr[1653] = 8'b00100000;
		color_arr[1654] = 8'b00100000;
		color_arr[1655] = 8'b00100000;
		color_arr[1656] = 8'b00100000;
		color_arr[1657] = 8'b00100000;
		color_arr[1658] = 8'b00100000;
		color_arr[1659] = 8'b00100000;
		color_arr[1660] = 8'b00100000;
		color_arr[1661] = 8'b00100000;
		color_arr[1662] = 8'b00100000;
		color_arr[1663] = 8'b00100000;
		color_arr[1664] = 8'b00010010;
		color_arr[1665] = 8'b00010010;
		color_arr[1666] = 8'b00010010;
		color_arr[1667] = 8'b00010010;
		color_arr[1668] = 8'b00010010;
		color_arr[1669] = 8'b00010010;
		color_arr[1670] = 8'b00010010;
		color_arr[1671] = 8'b00010010;
		color_arr[1672] = 8'b00000010;
		color_arr[1673] = 8'b00000010;
		color_arr[1674] = 8'b00000010;
		color_arr[1675] = 8'b00000010;
		color_arr[1676] = 8'b00000010;
		color_arr[1677] = 8'b00000010;
		color_arr[1678] = 8'b00000010;
		color_arr[1679] = 8'b00000010;
		color_arr[1680] = 8'b00000010;
		color_arr[1681] = 8'b00000010;
		color_arr[1682] = 8'b00000010;
		color_arr[1683] = 8'b00000010;
		color_arr[1684] = 8'b00000010;
		color_arr[1685] = 8'b00000010;
		color_arr[1686] = 8'b00000010;
		color_arr[1687] = 8'b00000000;
		color_arr[1688] = 8'b00000000;
		color_arr[1689] = 8'b00000000;
		color_arr[1690] = 8'b00000000;
		color_arr[1691] = 8'b00000010;
		color_arr[1692] = 8'b00000010;
		color_arr[1693] = 8'b00000010;
		color_arr[1694] = 8'b00000010;
		color_arr[1695] = 8'b00000010;
		color_arr[1696] = 8'b00000010;
		color_arr[1697] = 8'b00000010;
		color_arr[1698] = 8'b00000010;
		color_arr[1699] = 8'b00000010;
		color_arr[1700] = 8'b00000010;
		color_arr[1701] = 8'b00000010;
		color_arr[1702] = 8'b00100000;
		color_arr[1703] = 8'b00100000;
		color_arr[1704] = 8'b00100000;
		color_arr[1705] = 8'b00100000;
		color_arr[1706] = 8'b00100000;
		color_arr[1707] = 8'b00100000;
		color_arr[1708] = 8'b00100000;
		color_arr[1709] = 8'b00100000;
		color_arr[1710] = 8'b00100000;
		color_arr[1711] = 8'b00100000;
		color_arr[1712] = 8'b00100000;
		color_arr[1713] = 8'b00100000;
		color_arr[1714] = 8'b00100000;
		color_arr[1715] = 8'b00100000;
		color_arr[1716] = 8'b00100000;
		color_arr[1717] = 8'b00100000;
		color_arr[1718] = 8'b00100000;
		color_arr[1719] = 8'b00100000;
		color_arr[1720] = 8'b00100000;
		color_arr[1721] = 8'b00100000;
		color_arr[1722] = 8'b00100000;
		color_arr[1723] = 8'b00100000;
		color_arr[1724] = 8'b00100000;
		color_arr[1725] = 8'b00100000;
		color_arr[1726] = 8'b00100000;
		color_arr[1727] = 8'b00100000;
		color_arr[1728] = 8'b00010010;
		color_arr[1729] = 8'b00010010;
		color_arr[1730] = 8'b00010010;
		color_arr[1731] = 8'b00010010;
		color_arr[1732] = 8'b00010010;
		color_arr[1733] = 8'b00010010;
		color_arr[1734] = 8'b00010010;
		color_arr[1735] = 8'b00010010;
		color_arr[1736] = 8'b00000010;
		color_arr[1737] = 8'b00000010;
		color_arr[1738] = 8'b00000010;
		color_arr[1739] = 8'b00000010;
		color_arr[1740] = 8'b00000010;
		color_arr[1741] = 8'b00000010;
		color_arr[1742] = 8'b00000010;
		color_arr[1743] = 8'b00000010;
		color_arr[1744] = 8'b00000010;
		color_arr[1745] = 8'b00000000;
		color_arr[1746] = 8'b00000000;
		color_arr[1747] = 8'b00000000;
		color_arr[1748] = 8'b00000000;
		color_arr[1749] = 8'b00000000;
		color_arr[1750] = 8'b00000000;
		color_arr[1751] = 8'b00000000;
		color_arr[1752] = 8'b00000000;
		color_arr[1753] = 8'b00000000;
		color_arr[1754] = 8'b00000010;
		color_arr[1755] = 8'b00000010;
		color_arr[1756] = 8'b00000010;
		color_arr[1757] = 8'b00000010;
		color_arr[1758] = 8'b00000010;
		color_arr[1759] = 8'b00000010;
		color_arr[1760] = 8'b00000010;
		color_arr[1761] = 8'b00000010;
		color_arr[1762] = 8'b00000010;
		color_arr[1763] = 8'b00000010;
		color_arr[1764] = 8'b00000010;
		color_arr[1765] = 8'b00000010;
		color_arr[1766] = 8'b00100000;
		color_arr[1767] = 8'b00100000;
		color_arr[1768] = 8'b00100000;
		color_arr[1769] = 8'b00100000;
		color_arr[1770] = 8'b00100000;
		color_arr[1771] = 8'b00100000;
		color_arr[1772] = 8'b00100000;
		color_arr[1773] = 8'b00100000;
		color_arr[1774] = 8'b00100000;
		color_arr[1775] = 8'b00100000;
		color_arr[1776] = 8'b00100000;
		color_arr[1777] = 8'b00100000;
		color_arr[1778] = 8'b00100000;
		color_arr[1779] = 8'b00100000;
		color_arr[1780] = 8'b00100000;
		color_arr[1781] = 8'b00100000;
		color_arr[1782] = 8'b00100000;
		color_arr[1783] = 8'b00100000;
		color_arr[1784] = 8'b00100000;
		color_arr[1785] = 8'b00100000;
		color_arr[1786] = 8'b00100000;
		color_arr[1787] = 8'b00100000;
		color_arr[1788] = 8'b00100000;
		color_arr[1789] = 8'b00100000;
		color_arr[1790] = 8'b00100000;
		color_arr[1791] = 8'b00100000;
		color_arr[1792] = 8'b00010010;
		color_arr[1793] = 8'b00010010;
		color_arr[1794] = 8'b00010010;
		color_arr[1795] = 8'b00010010;
		color_arr[1796] = 8'b00010010;
		color_arr[1797] = 8'b00010010;
		color_arr[1798] = 8'b00010010;
		color_arr[1799] = 8'b00010010;
		color_arr[1800] = 8'b00000010;
		color_arr[1801] = 8'b00000010;
		color_arr[1802] = 8'b00000010;
		color_arr[1803] = 8'b00000010;
		color_arr[1804] = 8'b00000010;
		color_arr[1805] = 8'b00000010;
		color_arr[1806] = 8'b00000010;
		color_arr[1807] = 8'b00000000;
		color_arr[1808] = 8'b00000000;
		color_arr[1809] = 8'b00000000;
		color_arr[1810] = 8'b00000000;
		color_arr[1811] = 8'b00000000;
		color_arr[1812] = 8'b00000000;
		color_arr[1813] = 8'b00000000;
		color_arr[1814] = 8'b00000000;
		color_arr[1815] = 8'b00000000;
		color_arr[1816] = 8'b00000010;
		color_arr[1817] = 8'b00000010;
		color_arr[1818] = 8'b00000010;
		color_arr[1819] = 8'b00000010;
		color_arr[1820] = 8'b00000010;
		color_arr[1821] = 8'b00000010;
		color_arr[1822] = 8'b00000010;
		color_arr[1823] = 8'b00000010;
		color_arr[1824] = 8'b00000010;
		color_arr[1825] = 8'b00000010;
		color_arr[1826] = 8'b00000010;
		color_arr[1827] = 8'b00000010;
		color_arr[1828] = 8'b00000010;
		color_arr[1829] = 8'b00000010;
		color_arr[1830] = 8'b00100000;
		color_arr[1831] = 8'b00100000;
		color_arr[1832] = 8'b00100000;
		color_arr[1833] = 8'b00100000;
		color_arr[1834] = 8'b00100000;
		color_arr[1835] = 8'b00100000;
		color_arr[1836] = 8'b00100000;
		color_arr[1837] = 8'b00100000;
		color_arr[1838] = 8'b00100000;
		color_arr[1839] = 8'b00100000;
		color_arr[1840] = 8'b00100000;
		color_arr[1841] = 8'b00100000;
		color_arr[1842] = 8'b00100000;
		color_arr[1843] = 8'b00100000;
		color_arr[1844] = 8'b00100000;
		color_arr[1845] = 8'b00100000;
		color_arr[1846] = 8'b00100000;
		color_arr[1847] = 8'b00100000;
		color_arr[1848] = 8'b00100000;
		color_arr[1849] = 8'b00100000;
		color_arr[1850] = 8'b00100000;
		color_arr[1851] = 8'b00100000;
		color_arr[1852] = 8'b00100000;
		color_arr[1853] = 8'b00100000;
		color_arr[1854] = 8'b00100000;
		color_arr[1855] = 8'b00100000;
		color_arr[1856] = 8'b00010010;
		color_arr[1857] = 8'b00010010;
		color_arr[1858] = 8'b00010010;
		color_arr[1859] = 8'b00010010;
		color_arr[1860] = 8'b00010010;
		color_arr[1861] = 8'b00010010;
		color_arr[1862] = 8'b00010010;
		color_arr[1863] = 8'b00010010;
		color_arr[1864] = 8'b00000010;
		color_arr[1865] = 8'b00000010;
		color_arr[1866] = 8'b00000010;
		color_arr[1867] = 8'b00000010;
		color_arr[1868] = 8'b00000010;
		color_arr[1869] = 8'b00000000;
		color_arr[1870] = 8'b00000000;
		color_arr[1871] = 8'b00000000;
		color_arr[1872] = 8'b00000000;
		color_arr[1873] = 8'b00000000;
		color_arr[1874] = 8'b00000010;
		color_arr[1875] = 8'b00000010;
		color_arr[1876] = 8'b00000010;
		color_arr[1877] = 8'b00000000;
		color_arr[1878] = 8'b00000000;
		color_arr[1879] = 8'b00000010;
		color_arr[1880] = 8'b00000010;
		color_arr[1881] = 8'b00000010;
		color_arr[1882] = 8'b00000010;
		color_arr[1883] = 8'b00000010;
		color_arr[1884] = 8'b00000010;
		color_arr[1885] = 8'b00000010;
		color_arr[1886] = 8'b00000010;
		color_arr[1887] = 8'b00000010;
		color_arr[1888] = 8'b00000010;
		color_arr[1889] = 8'b00000010;
		color_arr[1890] = 8'b00000010;
		color_arr[1891] = 8'b00000010;
		color_arr[1892] = 8'b00000010;
		color_arr[1893] = 8'b00000010;
		color_arr[1894] = 8'b00100000;
		color_arr[1895] = 8'b00100000;
		color_arr[1896] = 8'b00100000;
		color_arr[1897] = 8'b00100000;
		color_arr[1898] = 8'b00100000;
		color_arr[1899] = 8'b00100000;
		color_arr[1900] = 8'b00100000;
		color_arr[1901] = 8'b00100000;
		color_arr[1902] = 8'b00100000;
		color_arr[1903] = 8'b00100000;
		color_arr[1904] = 8'b00100000;
		color_arr[1905] = 8'b00100000;
		color_arr[1906] = 8'b00100000;
		color_arr[1907] = 8'b00100000;
		color_arr[1908] = 8'b00100000;
		color_arr[1909] = 8'b00100000;
		color_arr[1910] = 8'b00100000;
		color_arr[1911] = 8'b00100000;
		color_arr[1912] = 8'b00100000;
		color_arr[1913] = 8'b00100000;
		color_arr[1914] = 8'b00100000;
		color_arr[1915] = 8'b00100000;
		color_arr[1916] = 8'b00100000;
		color_arr[1917] = 8'b00100000;
		color_arr[1918] = 8'b00100000;
		color_arr[1919] = 8'b00100000;
		color_arr[1920] = 8'b00010010;
		color_arr[1921] = 8'b00010010;
		color_arr[1922] = 8'b00010010;
		color_arr[1923] = 8'b00010010;
		color_arr[1924] = 8'b00010010;
		color_arr[1925] = 8'b00010010;
		color_arr[1926] = 8'b00010010;
		color_arr[1927] = 8'b00010010;
		color_arr[1928] = 8'b00000010;
		color_arr[1929] = 8'b00000010;
		color_arr[1930] = 8'b00000010;
		color_arr[1931] = 8'b00000010;
		color_arr[1932] = 8'b00000000;
		color_arr[1933] = 8'b00000000;
		color_arr[1934] = 8'b00000000;
		color_arr[1935] = 8'b00000000;
		color_arr[1936] = 8'b00000010;
		color_arr[1937] = 8'b00000010;
		color_arr[1938] = 8'b00000010;
		color_arr[1939] = 8'b00000010;
		color_arr[1940] = 8'b00000010;
		color_arr[1941] = 8'b00000010;
		color_arr[1942] = 8'b00000010;
		color_arr[1943] = 8'b00000010;
		color_arr[1944] = 8'b00000010;
		color_arr[1945] = 8'b00000010;
		color_arr[1946] = 8'b00000010;
		color_arr[1947] = 8'b00000010;
		color_arr[1948] = 8'b00000010;
		color_arr[1949] = 8'b00000010;
		color_arr[1950] = 8'b00000010;
		color_arr[1951] = 8'b00000010;
		color_arr[1952] = 8'b00000010;
		color_arr[1953] = 8'b00000010;
		color_arr[1954] = 8'b00000010;
		color_arr[1955] = 8'b00000010;
		color_arr[1956] = 8'b00000010;
		color_arr[1957] = 8'b00000010;
		color_arr[1958] = 8'b00100000;
		color_arr[1959] = 8'b00100000;
		color_arr[1960] = 8'b00100000;
		color_arr[1961] = 8'b00100000;
		color_arr[1962] = 8'b00100000;
		color_arr[1963] = 8'b00100000;
		color_arr[1964] = 8'b00100000;
		color_arr[1965] = 8'b00100000;
		color_arr[1966] = 8'b00100000;
		color_arr[1967] = 8'b00100000;
		color_arr[1968] = 8'b00100000;
		color_arr[1969] = 8'b00100000;
		color_arr[1970] = 8'b00100000;
		color_arr[1971] = 8'b00100000;
		color_arr[1972] = 8'b00100000;
		color_arr[1973] = 8'b00100000;
		color_arr[1974] = 8'b00100000;
		color_arr[1975] = 8'b00100000;
		color_arr[1976] = 8'b00100000;
		color_arr[1977] = 8'b00100000;
		color_arr[1978] = 8'b00100000;
		color_arr[1979] = 8'b00100000;
		color_arr[1980] = 8'b00100000;
		color_arr[1981] = 8'b00100000;
		color_arr[1982] = 8'b00100000;
		color_arr[1983] = 8'b00100000;
		color_arr[1984] = 8'b00010010;
		color_arr[1985] = 8'b00010010;
		color_arr[1986] = 8'b00010010;
		color_arr[1987] = 8'b00010010;
		color_arr[1988] = 8'b00010010;
		color_arr[1989] = 8'b00010010;
		color_arr[1990] = 8'b00010010;
		color_arr[1991] = 8'b00010010;
		color_arr[1992] = 8'b00000010;
		color_arr[1993] = 8'b00000010;
		color_arr[1994] = 8'b00000000;
		color_arr[1995] = 8'b00000000;
		color_arr[1996] = 8'b00000000;
		color_arr[1997] = 8'b00000000;
		color_arr[1998] = 8'b00000010;
		color_arr[1999] = 8'b00000010;
		color_arr[2000] = 8'b00000010;
		color_arr[2001] = 8'b00000010;
		color_arr[2002] = 8'b00000010;
		color_arr[2003] = 8'b00000010;
		color_arr[2004] = 8'b00000010;
		color_arr[2005] = 8'b00000010;
		color_arr[2006] = 8'b00000010;
		color_arr[2007] = 8'b00000010;
		color_arr[2008] = 8'b00000010;
		color_arr[2009] = 8'b00000010;
		color_arr[2010] = 8'b00000010;
		color_arr[2011] = 8'b00000010;
		color_arr[2012] = 8'b00000010;
		color_arr[2013] = 8'b00000010;
		color_arr[2014] = 8'b00000010;
		color_arr[2015] = 8'b00000010;
		color_arr[2016] = 8'b00000010;
		color_arr[2017] = 8'b00000010;
		color_arr[2018] = 8'b00000010;
		color_arr[2019] = 8'b00000010;
		color_arr[2020] = 8'b00000010;
		color_arr[2021] = 8'b00000010;
		color_arr[2022] = 8'b00100000;
		color_arr[2023] = 8'b00100000;
		color_arr[2024] = 8'b00100000;
		color_arr[2025] = 8'b00100000;
		color_arr[2026] = 8'b00100000;
		color_arr[2027] = 8'b00100000;
		color_arr[2028] = 8'b00100000;
		color_arr[2029] = 8'b00100000;
		color_arr[2030] = 8'b00100000;
		color_arr[2031] = 8'b00100000;
		color_arr[2032] = 8'b00100000;
		color_arr[2033] = 8'b00100000;
		color_arr[2034] = 8'b00100000;
		color_arr[2035] = 8'b00100000;
		color_arr[2036] = 8'b00100000;
		color_arr[2037] = 8'b00100000;
		color_arr[2038] = 8'b00000000;
		color_arr[2039] = 8'b00000000;
		color_arr[2040] = 8'b00000000;
		color_arr[2041] = 8'b00000000;
		color_arr[2042] = 8'b00000000;
		color_arr[2043] = 8'b00000000;
		color_arr[2044] = 8'b00000000;
		color_arr[2045] = 8'b00000000;
		color_arr[2046] = 8'b00000000;
		color_arr[2047] = 8'b00000000;
		color_arr[2048] = 8'b00010010;
		color_arr[2049] = 8'b00010010;
		color_arr[2050] = 8'b00010010;
		color_arr[2051] = 8'b00010010;
		color_arr[2052] = 8'b00010010;
		color_arr[2053] = 8'b00010010;
		color_arr[2054] = 8'b00010010;
		color_arr[2055] = 8'b00010010;
		color_arr[2056] = 8'b00000010;
		color_arr[2057] = 8'b00000000;
		color_arr[2058] = 8'b00000000;
		color_arr[2059] = 8'b00000000;
		color_arr[2060] = 8'b00000000;
		color_arr[2061] = 8'b00000010;
		color_arr[2062] = 8'b00000010;
		color_arr[2063] = 8'b00000010;
		color_arr[2064] = 8'b00000010;
		color_arr[2065] = 8'b00000010;
		color_arr[2066] = 8'b00000010;
		color_arr[2067] = 8'b00000010;
		color_arr[2068] = 8'b00000010;
		color_arr[2069] = 8'b00000010;
		color_arr[2070] = 8'b00000010;
		color_arr[2071] = 8'b00000010;
		color_arr[2072] = 8'b00000010;
		color_arr[2073] = 8'b00000010;
		color_arr[2074] = 8'b00000010;
		color_arr[2075] = 8'b00000010;
		color_arr[2076] = 8'b00000010;
		color_arr[2077] = 8'b00000010;
		color_arr[2078] = 8'b00000010;
		color_arr[2079] = 8'b00000010;
		color_arr[2080] = 8'b00000010;
		color_arr[2081] = 8'b00000010;
		color_arr[2082] = 8'b00000010;
		color_arr[2083] = 8'b00000010;
		color_arr[2084] = 8'b00000010;
		color_arr[2085] = 8'b00000010;
		color_arr[2086] = 8'b00100000;
		color_arr[2087] = 8'b00100000;
		color_arr[2088] = 8'b00100000;
		color_arr[2089] = 8'b00100000;
		color_arr[2090] = 8'b00100000;
		color_arr[2091] = 8'b00100000;
		color_arr[2092] = 8'b00100000;
		color_arr[2093] = 8'b00100000;
		color_arr[2094] = 8'b00100000;
		color_arr[2095] = 8'b00100000;
		color_arr[2096] = 8'b00000000;
		color_arr[2097] = 8'b00000000;
		color_arr[2098] = 8'b00000000;
		color_arr[2099] = 8'b00000000;
		color_arr[2100] = 8'b00000000;
		color_arr[2101] = 8'b00000000;
		color_arr[2102] = 8'b00000000;
		color_arr[2103] = 8'b00000000;
		color_arr[2104] = 8'b00000000;
		color_arr[2105] = 8'b00000000;
		color_arr[2106] = 8'b00000000;
		color_arr[2107] = 8'b00000000;
		color_arr[2108] = 8'b00000000;
		color_arr[2109] = 8'b00000000;
		color_arr[2110] = 8'b00000000;
		color_arr[2111] = 8'b00000000;
		color_arr[2112] = 8'b00010010;
		color_arr[2113] = 8'b00010010;
		color_arr[2114] = 8'b00010010;
		color_arr[2115] = 8'b00010010;
		color_arr[2116] = 8'b00010010;
		color_arr[2117] = 8'b00010010;
		color_arr[2118] = 8'b00010010;
		color_arr[2119] = 8'b00010010;
		color_arr[2120] = 8'b00000000;
		color_arr[2121] = 8'b00000000;
		color_arr[2122] = 8'b00000000;
		color_arr[2123] = 8'b00000010;
		color_arr[2124] = 8'b00000010;
		color_arr[2125] = 8'b00000010;
		color_arr[2126] = 8'b00000010;
		color_arr[2127] = 8'b00000010;
		color_arr[2128] = 8'b00000010;
		color_arr[2129] = 8'b00000010;
		color_arr[2130] = 8'b00000010;
		color_arr[2131] = 8'b00000010;
		color_arr[2132] = 8'b00000010;
		color_arr[2133] = 8'b00000010;
		color_arr[2134] = 8'b00000010;
		color_arr[2135] = 8'b00000010;
		color_arr[2136] = 8'b00000010;
		color_arr[2137] = 8'b00000010;
		color_arr[2138] = 8'b00000010;
		color_arr[2139] = 8'b00000010;
		color_arr[2140] = 8'b00000010;
		color_arr[2141] = 8'b00000010;
		color_arr[2142] = 8'b00000010;
		color_arr[2143] = 8'b00000010;
		color_arr[2144] = 8'b00000010;
		color_arr[2145] = 8'b00000010;
		color_arr[2146] = 8'b00000010;
		color_arr[2147] = 8'b00000010;
		color_arr[2148] = 8'b00000010;
		color_arr[2149] = 8'b00000010;
		color_arr[2150] = 8'b00100000;
		color_arr[2151] = 8'b00100000;
		color_arr[2152] = 8'b00100000;
		color_arr[2153] = 8'b00100000;
		color_arr[2154] = 8'b00100000;
		color_arr[2155] = 8'b00000000;
		color_arr[2156] = 8'b00000000;
		color_arr[2157] = 8'b00000000;
		color_arr[2158] = 8'b00000000;
		color_arr[2159] = 8'b00000000;
		color_arr[2160] = 8'b00000000;
		color_arr[2161] = 8'b00000000;
		color_arr[2162] = 8'b00000000;
		color_arr[2163] = 8'b00000000;
		color_arr[2164] = 8'b00000000;
		color_arr[2165] = 8'b00000000;
		color_arr[2166] = 8'b00000000;
		color_arr[2167] = 8'b00100000;
		color_arr[2168] = 8'b00100000;
		color_arr[2169] = 8'b00100000;
		color_arr[2170] = 8'b00100000;
		color_arr[2171] = 8'b00100000;
		color_arr[2172] = 8'b00100000;
		color_arr[2173] = 8'b00100000;
		color_arr[2174] = 8'b00100000;
		color_arr[2175] = 8'b00100000;
		color_arr[2176] = 8'b00010010;
		color_arr[2177] = 8'b00010010;
		color_arr[2178] = 8'b00010010;
		color_arr[2179] = 8'b00010010;
		color_arr[2180] = 8'b00010010;
		color_arr[2181] = 8'b00010010;
		color_arr[2182] = 8'b00010010;
		color_arr[2183] = 8'b00000000;
		color_arr[2184] = 8'b00000000;
		color_arr[2185] = 8'b00000000;
		color_arr[2186] = 8'b00000010;
		color_arr[2187] = 8'b00000010;
		color_arr[2188] = 8'b00000010;
		color_arr[2189] = 8'b00000010;
		color_arr[2190] = 8'b00000010;
		color_arr[2191] = 8'b00000010;
		color_arr[2192] = 8'b00000010;
		color_arr[2193] = 8'b00000010;
		color_arr[2194] = 8'b00000010;
		color_arr[2195] = 8'b00000010;
		color_arr[2196] = 8'b00000010;
		color_arr[2197] = 8'b00000010;
		color_arr[2198] = 8'b00000010;
		color_arr[2199] = 8'b00000010;
		color_arr[2200] = 8'b00000010;
		color_arr[2201] = 8'b00000010;
		color_arr[2202] = 8'b00000010;
		color_arr[2203] = 8'b00000010;
		color_arr[2204] = 8'b00000010;
		color_arr[2205] = 8'b00000010;
		color_arr[2206] = 8'b00000010;
		color_arr[2207] = 8'b00000010;
		color_arr[2208] = 8'b00000010;
		color_arr[2209] = 8'b00000010;
		color_arr[2210] = 8'b00000010;
		color_arr[2211] = 8'b00000010;
		color_arr[2212] = 8'b00000010;
		color_arr[2213] = 8'b00000010;
		color_arr[2214] = 8'b00100000;
		color_arr[2215] = 8'b00000000;
		color_arr[2216] = 8'b00000000;
		color_arr[2217] = 8'b00000000;
		color_arr[2218] = 8'b00000000;
		color_arr[2219] = 8'b00000000;
		color_arr[2220] = 8'b00000000;
		color_arr[2221] = 8'b00000000;
		color_arr[2222] = 8'b00000000;
		color_arr[2223] = 8'b00000000;
		color_arr[2224] = 8'b00000000;
		color_arr[2225] = 8'b00100000;
		color_arr[2226] = 8'b00100000;
		color_arr[2227] = 8'b00100000;
		color_arr[2228] = 8'b00100000;
		color_arr[2229] = 8'b00100000;
		color_arr[2230] = 8'b00100000;
		color_arr[2231] = 8'b00100000;
		color_arr[2232] = 8'b00100000;
		color_arr[2233] = 8'b00100000;
		color_arr[2234] = 8'b00100000;
		color_arr[2235] = 8'b00100000;
		color_arr[2236] = 8'b00100000;
		color_arr[2237] = 8'b00100000;
		color_arr[2238] = 8'b00100000;
		color_arr[2239] = 8'b00100000;
		color_arr[2240] = 8'b00010010;
		color_arr[2241] = 8'b00010010;
		color_arr[2242] = 8'b00010010;
		color_arr[2243] = 8'b00010010;
		color_arr[2244] = 8'b00010010;
		color_arr[2245] = 8'b00010010;
		color_arr[2246] = 8'b00000000;
		color_arr[2247] = 8'b00000000;
		color_arr[2248] = 8'b00000000;
		color_arr[2249] = 8'b00000010;
		color_arr[2250] = 8'b00000010;
		color_arr[2251] = 8'b00000010;
		color_arr[2252] = 8'b00000010;
		color_arr[2253] = 8'b00000010;
		color_arr[2254] = 8'b00000010;
		color_arr[2255] = 8'b00000010;
		color_arr[2256] = 8'b00000010;
		color_arr[2257] = 8'b00000010;
		color_arr[2258] = 8'b00000010;
		color_arr[2259] = 8'b00000010;
		color_arr[2260] = 8'b00000010;
		color_arr[2261] = 8'b00000010;
		color_arr[2262] = 8'b00000010;
		color_arr[2263] = 8'b00000010;
		color_arr[2264] = 8'b00000010;
		color_arr[2265] = 8'b00000010;
		color_arr[2266] = 8'b00000010;
		color_arr[2267] = 8'b00000010;
		color_arr[2268] = 8'b00000010;
		color_arr[2269] = 8'b00000010;
		color_arr[2270] = 8'b00000010;
		color_arr[2271] = 8'b00000010;
		color_arr[2272] = 8'b00000010;
		color_arr[2273] = 8'b00000010;
		color_arr[2274] = 8'b00000010;
		color_arr[2275] = 8'b00000010;
		color_arr[2276] = 8'b00000000;
		color_arr[2277] = 8'b00000000;
		color_arr[2278] = 8'b00000000;
		color_arr[2279] = 8'b00000000;
		color_arr[2280] = 8'b00000000;
		color_arr[2281] = 8'b00000000;
		color_arr[2282] = 8'b00000000;
		color_arr[2283] = 8'b00000000;
		color_arr[2284] = 8'b00100000;
		color_arr[2285] = 8'b00100000;
		color_arr[2286] = 8'b00100000;
		color_arr[2287] = 8'b00100000;
		color_arr[2288] = 8'b00100000;
		color_arr[2289] = 8'b00100000;
		color_arr[2290] = 8'b00100000;
		color_arr[2291] = 8'b00100000;
		color_arr[2292] = 8'b00100000;
		color_arr[2293] = 8'b00100000;
		color_arr[2294] = 8'b00100000;
		color_arr[2295] = 8'b00100000;
		color_arr[2296] = 8'b00100000;
		color_arr[2297] = 8'b00100000;
		color_arr[2298] = 8'b00100000;
		color_arr[2299] = 8'b00100000;
		color_arr[2300] = 8'b00100000;
		color_arr[2301] = 8'b00100000;
		color_arr[2302] = 8'b00100000;
		color_arr[2303] = 8'b00100000;
		color_arr[2304] = 8'b00010010;
		color_arr[2305] = 8'b00010010;
		color_arr[2306] = 8'b00010010;
		color_arr[2307] = 8'b00010010;
		color_arr[2308] = 8'b00010010;
		color_arr[2309] = 8'b00000000;
		color_arr[2310] = 8'b00000000;
		color_arr[2311] = 8'b00000000;
		color_arr[2312] = 8'b00000010;
		color_arr[2313] = 8'b00000010;
		color_arr[2314] = 8'b00000010;
		color_arr[2315] = 8'b00000010;
		color_arr[2316] = 8'b00000010;
		color_arr[2317] = 8'b00000010;
		color_arr[2318] = 8'b00000010;
		color_arr[2319] = 8'b00000010;
		color_arr[2320] = 8'b00000010;
		color_arr[2321] = 8'b00000010;
		color_arr[2322] = 8'b00000010;
		color_arr[2323] = 8'b00000010;
		color_arr[2324] = 8'b00000010;
		color_arr[2325] = 8'b00000010;
		color_arr[2326] = 8'b00000010;
		color_arr[2327] = 8'b00000010;
		color_arr[2328] = 8'b00000010;
		color_arr[2329] = 8'b00000010;
		color_arr[2330] = 8'b00000010;
		color_arr[2331] = 8'b00000010;
		color_arr[2332] = 8'b00000010;
		color_arr[2333] = 8'b00000010;
		color_arr[2334] = 8'b00000010;
		color_arr[2335] = 8'b00000010;
		color_arr[2336] = 8'b00000010;
		color_arr[2337] = 8'b00000010;
		color_arr[2338] = 8'b00000000;
		color_arr[2339] = 8'b00000000;
		color_arr[2340] = 8'b00000000;
		color_arr[2341] = 8'b00000000;
		color_arr[2342] = 8'b00000000;
		color_arr[2343] = 8'b00000000;
		color_arr[2344] = 8'b00100000;
		color_arr[2345] = 8'b00100000;
		color_arr[2346] = 8'b00100000;
		color_arr[2347] = 8'b00100000;
		color_arr[2348] = 8'b00100000;
		color_arr[2349] = 8'b00100000;
		color_arr[2350] = 8'b00100000;
		color_arr[2351] = 8'b00100000;
		color_arr[2352] = 8'b00100000;
		color_arr[2353] = 8'b00100000;
		color_arr[2354] = 8'b00100000;
		color_arr[2355] = 8'b00100000;
		color_arr[2356] = 8'b00100000;
		color_arr[2357] = 8'b00100000;
		color_arr[2358] = 8'b00100000;
		color_arr[2359] = 8'b00100000;
		color_arr[2360] = 8'b00100000;
		color_arr[2361] = 8'b00100000;
		color_arr[2362] = 8'b00100000;
		color_arr[2363] = 8'b00100000;
		color_arr[2364] = 8'b00100000;
		color_arr[2365] = 8'b00100000;
		color_arr[2366] = 8'b00100000;
		color_arr[2367] = 8'b00100000;
		color_arr[2368] = 8'b00010010;
		color_arr[2369] = 8'b00010010;
		color_arr[2370] = 8'b00010010;
		color_arr[2371] = 8'b00010010;
		color_arr[2372] = 8'b00010010;
		color_arr[2373] = 8'b00000000;
		color_arr[2374] = 8'b00000000;
		color_arr[2375] = 8'b00010010;
		color_arr[2376] = 8'b00000010;
		color_arr[2377] = 8'b00000010;
		color_arr[2378] = 8'b00000010;
		color_arr[2379] = 8'b00000010;
		color_arr[2380] = 8'b00000010;
		color_arr[2381] = 8'b00000010;
		color_arr[2382] = 8'b00000010;
		color_arr[2383] = 8'b00000010;
		color_arr[2384] = 8'b00000010;
		color_arr[2385] = 8'b00000010;
		color_arr[2386] = 8'b00000010;
		color_arr[2387] = 8'b00000010;
		color_arr[2388] = 8'b00000010;
		color_arr[2389] = 8'b00000010;
		color_arr[2390] = 8'b00000010;
		color_arr[2391] = 8'b00000010;
		color_arr[2392] = 8'b00000010;
		color_arr[2393] = 8'b00000010;
		color_arr[2394] = 8'b00000010;
		color_arr[2395] = 8'b00000010;
		color_arr[2396] = 8'b00000010;
		color_arr[2397] = 8'b00000010;
		color_arr[2398] = 8'b00000010;
		color_arr[2399] = 8'b00000010;
		color_arr[2400] = 8'b00000000;
		color_arr[2401] = 8'b00000000;
		color_arr[2402] = 8'b00000000;
		color_arr[2403] = 8'b00000000;
		color_arr[2404] = 8'b00000000;
		color_arr[2405] = 8'b00000010;
		color_arr[2406] = 8'b00100000;
		color_arr[2407] = 8'b00100000;
		color_arr[2408] = 8'b00100000;
		color_arr[2409] = 8'b00100000;
		color_arr[2410] = 8'b00100000;
		color_arr[2411] = 8'b00100000;
		color_arr[2412] = 8'b00100000;
		color_arr[2413] = 8'b00100000;
		color_arr[2414] = 8'b00100000;
		color_arr[2415] = 8'b00100000;
		color_arr[2416] = 8'b00100000;
		color_arr[2417] = 8'b00100000;
		color_arr[2418] = 8'b00100000;
		color_arr[2419] = 8'b00100000;
		color_arr[2420] = 8'b00100000;
		color_arr[2421] = 8'b00100000;
		color_arr[2422] = 8'b00100000;
		color_arr[2423] = 8'b00100000;
		color_arr[2424] = 8'b00100000;
		color_arr[2425] = 8'b00100000;
		color_arr[2426] = 8'b00100000;
		color_arr[2427] = 8'b00100000;
		color_arr[2428] = 8'b00100000;
		color_arr[2429] = 8'b00100000;
		color_arr[2430] = 8'b00100000;
		color_arr[2431] = 8'b00100000;
		color_arr[2432] = 8'b00010010;
		color_arr[2433] = 8'b00010010;
		color_arr[2434] = 8'b00010010;
		color_arr[2435] = 8'b00010010;
		color_arr[2436] = 8'b00000000;
		color_arr[2437] = 8'b00000000;
		color_arr[2438] = 8'b00000000;
		color_arr[2439] = 8'b00010010;
		color_arr[2440] = 8'b00000010;
		color_arr[2441] = 8'b00000010;
		color_arr[2442] = 8'b00000010;
		color_arr[2443] = 8'b00000010;
		color_arr[2444] = 8'b00000010;
		color_arr[2445] = 8'b00000010;
		color_arr[2446] = 8'b00000010;
		color_arr[2447] = 8'b00000010;
		color_arr[2448] = 8'b00000010;
		color_arr[2449] = 8'b00000010;
		color_arr[2450] = 8'b00000010;
		color_arr[2451] = 8'b00000010;
		color_arr[2452] = 8'b00000010;
		color_arr[2453] = 8'b00000010;
		color_arr[2454] = 8'b00000010;
		color_arr[2455] = 8'b00000010;
		color_arr[2456] = 8'b00000010;
		color_arr[2457] = 8'b00000010;
		color_arr[2458] = 8'b00000010;
		color_arr[2459] = 8'b00000010;
		color_arr[2460] = 8'b00000010;
		color_arr[2461] = 8'b00000010;
		color_arr[2462] = 8'b00000010;
		color_arr[2463] = 8'b00000000;
		color_arr[2464] = 8'b00000000;
		color_arr[2465] = 8'b00000000;
		color_arr[2466] = 8'b00000000;
		color_arr[2467] = 8'b00000010;
		color_arr[2468] = 8'b00000010;
		color_arr[2469] = 8'b00000010;
		color_arr[2470] = 8'b00100000;
		color_arr[2471] = 8'b00100000;
		color_arr[2472] = 8'b00100000;
		color_arr[2473] = 8'b00100000;
		color_arr[2474] = 8'b00100000;
		color_arr[2475] = 8'b00100000;
		color_arr[2476] = 8'b00100000;
		color_arr[2477] = 8'b00100000;
		color_arr[2478] = 8'b00100000;
		color_arr[2479] = 8'b00100000;
		color_arr[2480] = 8'b00100000;
		color_arr[2481] = 8'b00100000;
		color_arr[2482] = 8'b00100000;
		color_arr[2483] = 8'b00100000;
		color_arr[2484] = 8'b00100000;
		color_arr[2485] = 8'b00100000;
		color_arr[2486] = 8'b00100000;
		color_arr[2487] = 8'b00100000;
		color_arr[2488] = 8'b00100000;
		color_arr[2489] = 8'b00100000;
		color_arr[2490] = 8'b00100000;
		color_arr[2491] = 8'b00100000;
		color_arr[2492] = 8'b00100000;
		color_arr[2493] = 8'b00100000;
		color_arr[2494] = 8'b00100000;
		color_arr[2495] = 8'b00100000;
		color_arr[2496] = 8'b00010010;
		color_arr[2497] = 8'b00010010;
		color_arr[2498] = 8'b00010010;
		color_arr[2499] = 8'b00010010;
		color_arr[2500] = 8'b00000000;
		color_arr[2501] = 8'b00000000;
		color_arr[2502] = 8'b00010010;
		color_arr[2503] = 8'b00010010;
		color_arr[2504] = 8'b00000010;
		color_arr[2505] = 8'b00000010;
		color_arr[2506] = 8'b00000010;
		color_arr[2507] = 8'b00000010;
		color_arr[2508] = 8'b00000010;
		color_arr[2509] = 8'b00000010;
		color_arr[2510] = 8'b00000010;
		color_arr[2511] = 8'b00000010;
		color_arr[2512] = 8'b00000010;
		color_arr[2513] = 8'b00000010;
		color_arr[2514] = 8'b00000010;
		color_arr[2515] = 8'b00000010;
		color_arr[2516] = 8'b00000010;
		color_arr[2517] = 8'b00000010;
		color_arr[2518] = 8'b00000010;
		color_arr[2519] = 8'b00000010;
		color_arr[2520] = 8'b00000010;
		color_arr[2521] = 8'b00000010;
		color_arr[2522] = 8'b00000010;
		color_arr[2523] = 8'b00000010;
		color_arr[2524] = 8'b00000010;
		color_arr[2525] = 8'b00000010;
		color_arr[2526] = 8'b00000000;
		color_arr[2527] = 8'b00000000;
		color_arr[2528] = 8'b00000000;
		color_arr[2529] = 8'b00000010;
		color_arr[2530] = 8'b00000010;
		color_arr[2531] = 8'b00000010;
		color_arr[2532] = 8'b00000010;
		color_arr[2533] = 8'b00000010;
		color_arr[2534] = 8'b00100000;
		color_arr[2535] = 8'b00100000;
		color_arr[2536] = 8'b00100000;
		color_arr[2537] = 8'b00100000;
		color_arr[2538] = 8'b00100000;
		color_arr[2539] = 8'b00100000;
		color_arr[2540] = 8'b00100000;
		color_arr[2541] = 8'b00100000;
		color_arr[2542] = 8'b00100000;
		color_arr[2543] = 8'b00100000;
		color_arr[2544] = 8'b00100000;
		color_arr[2545] = 8'b00100000;
		color_arr[2546] = 8'b00100000;
		color_arr[2547] = 8'b00100000;
		color_arr[2548] = 8'b00100000;
		color_arr[2549] = 8'b00100000;
		color_arr[2550] = 8'b00100000;
		color_arr[2551] = 8'b00100000;
		color_arr[2552] = 8'b00100000;
		color_arr[2553] = 8'b00100000;
		color_arr[2554] = 8'b00100000;
		color_arr[2555] = 8'b00100000;
		color_arr[2556] = 8'b00100000;
		color_arr[2557] = 8'b00100000;
		color_arr[2558] = 8'b00100000;
		color_arr[2559] = 8'b00100000;
		color_arr[2560] = 8'b00010010;
		color_arr[2561] = 8'b00010010;
		color_arr[2562] = 8'b00010010;
		color_arr[2563] = 8'b00000000;
		color_arr[2564] = 8'b00000000;
		color_arr[2565] = 8'b00000000;
		color_arr[2566] = 8'b00010010;
		color_arr[2567] = 8'b00010010;
		color_arr[2568] = 8'b00000010;
		color_arr[2569] = 8'b00000010;
		color_arr[2570] = 8'b00000010;
		color_arr[2571] = 8'b00000010;
		color_arr[2572] = 8'b00000010;
		color_arr[2573] = 8'b00000010;
		color_arr[2574] = 8'b00000010;
		color_arr[2575] = 8'b00000010;
		color_arr[2576] = 8'b00000010;
		color_arr[2577] = 8'b00000010;
		color_arr[2578] = 8'b00000010;
		color_arr[2579] = 8'b00000010;
		color_arr[2580] = 8'b00000010;
		color_arr[2581] = 8'b00000010;
		color_arr[2582] = 8'b00000010;
		color_arr[2583] = 8'b00000010;
		color_arr[2584] = 8'b00000010;
		color_arr[2585] = 8'b00000010;
		color_arr[2586] = 8'b00000010;
		color_arr[2587] = 8'b00000010;
		color_arr[2588] = 8'b00000000;
		color_arr[2589] = 8'b00000000;
		color_arr[2590] = 8'b00000000;
		color_arr[2591] = 8'b00000000;
		color_arr[2592] = 8'b00000010;
		color_arr[2593] = 8'b00000010;
		color_arr[2594] = 8'b00000010;
		color_arr[2595] = 8'b00000010;
		color_arr[2596] = 8'b00000010;
		color_arr[2597] = 8'b00000010;
		color_arr[2598] = 8'b00100000;
		color_arr[2599] = 8'b00100000;
		color_arr[2600] = 8'b00100000;
		color_arr[2601] = 8'b00100000;
		color_arr[2602] = 8'b00100000;
		color_arr[2603] = 8'b00100000;
		color_arr[2604] = 8'b00100000;
		color_arr[2605] = 8'b00100000;
		color_arr[2606] = 8'b00100000;
		color_arr[2607] = 8'b00100000;
		color_arr[2608] = 8'b00100000;
		color_arr[2609] = 8'b00100000;
		color_arr[2610] = 8'b00100000;
		color_arr[2611] = 8'b00100000;
		color_arr[2612] = 8'b00100000;
		color_arr[2613] = 8'b00100000;
		color_arr[2614] = 8'b00100000;
		color_arr[2615] = 8'b00100000;
		color_arr[2616] = 8'b00100000;
		color_arr[2617] = 8'b00100000;
		color_arr[2618] = 8'b00100000;
		color_arr[2619] = 8'b00100000;
		color_arr[2620] = 8'b00100000;
		color_arr[2621] = 8'b00100000;
		color_arr[2622] = 8'b00100000;
		color_arr[2623] = 8'b00100000;
		color_arr[2624] = 8'b00010010;
		color_arr[2625] = 8'b00010010;
		color_arr[2626] = 8'b00010010;
		color_arr[2627] = 8'b00000000;
		color_arr[2628] = 8'b00000000;
		color_arr[2629] = 8'b00010010;
		color_arr[2630] = 8'b00010010;
		color_arr[2631] = 8'b00010010;
		color_arr[2632] = 8'b00000010;
		color_arr[2633] = 8'b00000010;
		color_arr[2634] = 8'b00000010;
		color_arr[2635] = 8'b00000010;
		color_arr[2636] = 8'b00000010;
		color_arr[2637] = 8'b00000010;
		color_arr[2638] = 8'b00000010;
		color_arr[2639] = 8'b00000010;
		color_arr[2640] = 8'b00000010;
		color_arr[2641] = 8'b00000010;
		color_arr[2642] = 8'b00000010;
		color_arr[2643] = 8'b00000010;
		color_arr[2644] = 8'b00000010;
		color_arr[2645] = 8'b00000010;
		color_arr[2646] = 8'b00000010;
		color_arr[2647] = 8'b00000010;
		color_arr[2648] = 8'b00000010;
		color_arr[2649] = 8'b00000010;
		color_arr[2650] = 8'b00000010;
		color_arr[2651] = 8'b00000000;
		color_arr[2652] = 8'b00000000;
		color_arr[2653] = 8'b00000000;
		color_arr[2654] = 8'b00000000;
		color_arr[2655] = 8'b00000010;
		color_arr[2656] = 8'b00000010;
		color_arr[2657] = 8'b00000010;
		color_arr[2658] = 8'b00000010;
		color_arr[2659] = 8'b00000010;
		color_arr[2660] = 8'b00000010;
		color_arr[2661] = 8'b00000010;
		color_arr[2662] = 8'b00100000;
		color_arr[2663] = 8'b00100000;
		color_arr[2664] = 8'b00100000;
		color_arr[2665] = 8'b00100000;
		color_arr[2666] = 8'b00100000;
		color_arr[2667] = 8'b00100000;
		color_arr[2668] = 8'b00100000;
		color_arr[2669] = 8'b00100000;
		color_arr[2670] = 8'b00100000;
		color_arr[2671] = 8'b00100000;
		color_arr[2672] = 8'b00100000;
		color_arr[2673] = 8'b00100000;
		color_arr[2674] = 8'b00100000;
		color_arr[2675] = 8'b00100000;
		color_arr[2676] = 8'b00100000;
		color_arr[2677] = 8'b00100000;
		color_arr[2678] = 8'b00100000;
		color_arr[2679] = 8'b00100000;
		color_arr[2680] = 8'b00100000;
		color_arr[2681] = 8'b00100000;
		color_arr[2682] = 8'b00100000;
		color_arr[2683] = 8'b00100000;
		color_arr[2684] = 8'b00100000;
		color_arr[2685] = 8'b00100000;
		color_arr[2686] = 8'b00100000;
		color_arr[2687] = 8'b00100000;
		color_arr[2688] = 8'b00010010;
		color_arr[2689] = 8'b00010010;
		color_arr[2690] = 8'b00010010;
		color_arr[2691] = 8'b00000000;
		color_arr[2692] = 8'b00000000;
		color_arr[2693] = 8'b00010010;
		color_arr[2694] = 8'b00010010;
		color_arr[2695] = 8'b00010010;
		color_arr[2696] = 8'b00000010;
		color_arr[2697] = 8'b00000010;
		color_arr[2698] = 8'b00000010;
		color_arr[2699] = 8'b00000010;
		color_arr[2700] = 8'b00000010;
		color_arr[2701] = 8'b00000010;
		color_arr[2702] = 8'b00000010;
		color_arr[2703] = 8'b00000010;
		color_arr[2704] = 8'b00000010;
		color_arr[2705] = 8'b00000010;
		color_arr[2706] = 8'b00000010;
		color_arr[2707] = 8'b00000010;
		color_arr[2708] = 8'b00000010;
		color_arr[2709] = 8'b00000010;
		color_arr[2710] = 8'b00000010;
		color_arr[2711] = 8'b00000010;
		color_arr[2712] = 8'b00000010;
		color_arr[2713] = 8'b00000010;
		color_arr[2714] = 8'b00000000;
		color_arr[2715] = 8'b00000000;
		color_arr[2716] = 8'b00000000;
		color_arr[2717] = 8'b00000010;
		color_arr[2718] = 8'b00000010;
		color_arr[2719] = 8'b00000010;
		color_arr[2720] = 8'b00000010;
		color_arr[2721] = 8'b00000010;
		color_arr[2722] = 8'b00000010;
		color_arr[2723] = 8'b00000010;
		color_arr[2724] = 8'b00000010;
		color_arr[2725] = 8'b00000010;
		color_arr[2726] = 8'b00100000;
		color_arr[2727] = 8'b00100000;
		color_arr[2728] = 8'b00100000;
		color_arr[2729] = 8'b00100000;
		color_arr[2730] = 8'b00100000;
		color_arr[2731] = 8'b00100000;
		color_arr[2732] = 8'b00100000;
		color_arr[2733] = 8'b00100000;
		color_arr[2734] = 8'b00100000;
		color_arr[2735] = 8'b00100000;
		color_arr[2736] = 8'b00100000;
		color_arr[2737] = 8'b00100000;
		color_arr[2738] = 8'b00100000;
		color_arr[2739] = 8'b00100000;
		color_arr[2740] = 8'b00100000;
		color_arr[2741] = 8'b00100000;
		color_arr[2742] = 8'b00100000;
		color_arr[2743] = 8'b00100000;
		color_arr[2744] = 8'b00100000;
		color_arr[2745] = 8'b00100000;
		color_arr[2746] = 8'b00100000;
		color_arr[2747] = 8'b00100000;
		color_arr[2748] = 8'b00100000;
		color_arr[2749] = 8'b00100000;
		color_arr[2750] = 8'b00100000;
		color_arr[2751] = 8'b00100000;
		color_arr[2752] = 8'b00010010;
		color_arr[2753] = 8'b00010010;
		color_arr[2754] = 8'b00010010;
		color_arr[2755] = 8'b00000000;
		color_arr[2756] = 8'b00000000;
		color_arr[2757] = 8'b00010010;
		color_arr[2758] = 8'b00010010;
		color_arr[2759] = 8'b00010010;
		color_arr[2760] = 8'b00000010;
		color_arr[2761] = 8'b00000010;
		color_arr[2762] = 8'b00000010;
		color_arr[2763] = 8'b00000010;
		color_arr[2764] = 8'b00000010;
		color_arr[2765] = 8'b00000010;
		color_arr[2766] = 8'b00000010;
		color_arr[2767] = 8'b00000010;
		color_arr[2768] = 8'b00000010;
		color_arr[2769] = 8'b00000010;
		color_arr[2770] = 8'b00000010;
		color_arr[2771] = 8'b00000010;
		color_arr[2772] = 8'b00000010;
		color_arr[2773] = 8'b00000010;
		color_arr[2774] = 8'b00000010;
		color_arr[2775] = 8'b00000010;
		color_arr[2776] = 8'b00000010;
		color_arr[2777] = 8'b00000010;
		color_arr[2778] = 8'b00000000;
		color_arr[2779] = 8'b00000000;
		color_arr[2780] = 8'b00000010;
		color_arr[2781] = 8'b00000010;
		color_arr[2782] = 8'b00000010;
		color_arr[2783] = 8'b00000010;
		color_arr[2784] = 8'b00000010;
		color_arr[2785] = 8'b00000010;
		color_arr[2786] = 8'b00000010;
		color_arr[2787] = 8'b00000010;
		color_arr[2788] = 8'b00000010;
		color_arr[2789] = 8'b00000010;
		color_arr[2790] = 8'b00100000;
		color_arr[2791] = 8'b00100000;
		color_arr[2792] = 8'b00100000;
		color_arr[2793] = 8'b00100000;
		color_arr[2794] = 8'b00100000;
		color_arr[2795] = 8'b00100000;
		color_arr[2796] = 8'b00100000;
		color_arr[2797] = 8'b00100000;
		color_arr[2798] = 8'b00100000;
		color_arr[2799] = 8'b00100000;
		color_arr[2800] = 8'b00100000;
		color_arr[2801] = 8'b00100000;
		color_arr[2802] = 8'b00100000;
		color_arr[2803] = 8'b00100000;
		color_arr[2804] = 8'b00100000;
		color_arr[2805] = 8'b00100000;
		color_arr[2806] = 8'b00100000;
		color_arr[2807] = 8'b00100000;
		color_arr[2808] = 8'b00100000;
		color_arr[2809] = 8'b00100000;
		color_arr[2810] = 8'b00100000;
		color_arr[2811] = 8'b00100000;
		color_arr[2812] = 8'b00100000;
		color_arr[2813] = 8'b00100000;
		color_arr[2814] = 8'b00100000;
		color_arr[2815] = 8'b00100000;
		color_arr[2816] = 8'b00010010;
		color_arr[2817] = 8'b00010010;
		color_arr[2818] = 8'b00000000;
		color_arr[2819] = 8'b00000000;
		color_arr[2820] = 8'b00000000;
		color_arr[2821] = 8'b00010010;
		color_arr[2822] = 8'b00010010;
		color_arr[2823] = 8'b00010010;
		color_arr[2824] = 8'b00000010;
		color_arr[2825] = 8'b00000010;
		color_arr[2826] = 8'b00000010;
		color_arr[2827] = 8'b00000010;
		color_arr[2828] = 8'b00000010;
		color_arr[2829] = 8'b00000010;
		color_arr[2830] = 8'b00000010;
		color_arr[2831] = 8'b00000010;
		color_arr[2832] = 8'b00000010;
		color_arr[2833] = 8'b00000010;
		color_arr[2834] = 8'b00000010;
		color_arr[2835] = 8'b00000010;
		color_arr[2836] = 8'b00000010;
		color_arr[2837] = 8'b00000010;
		color_arr[2838] = 8'b00000010;
		color_arr[2839] = 8'b00000010;
		color_arr[2840] = 8'b00000010;
		color_arr[2841] = 8'b00000000;
		color_arr[2842] = 8'b00000000;
		color_arr[2843] = 8'b00000000;
		color_arr[2844] = 8'b00000010;
		color_arr[2845] = 8'b00000010;
		color_arr[2846] = 8'b00000010;
		color_arr[2847] = 8'b00000010;
		color_arr[2848] = 8'b00000010;
		color_arr[2849] = 8'b00000010;
		color_arr[2850] = 8'b00000010;
		color_arr[2851] = 8'b00000010;
		color_arr[2852] = 8'b00000010;
		color_arr[2853] = 8'b00000010;
		color_arr[2854] = 8'b00100000;
		color_arr[2855] = 8'b00100000;
		color_arr[2856] = 8'b00100000;
		color_arr[2857] = 8'b00100000;
		color_arr[2858] = 8'b00100000;
		color_arr[2859] = 8'b00100000;
		color_arr[2860] = 8'b00100000;
		color_arr[2861] = 8'b00100000;
		color_arr[2862] = 8'b00100000;
		color_arr[2863] = 8'b00100000;
		color_arr[2864] = 8'b00100000;
		color_arr[2865] = 8'b00100000;
		color_arr[2866] = 8'b00100000;
		color_arr[2867] = 8'b00100000;
		color_arr[2868] = 8'b00100000;
		color_arr[2869] = 8'b00100000;
		color_arr[2870] = 8'b00100000;
		color_arr[2871] = 8'b00100000;
		color_arr[2872] = 8'b00100000;
		color_arr[2873] = 8'b00100000;
		color_arr[2874] = 8'b00100000;
		color_arr[2875] = 8'b00100000;
		color_arr[2876] = 8'b00100000;
		color_arr[2877] = 8'b00100000;
		color_arr[2878] = 8'b00100000;
		color_arr[2879] = 8'b00100000;
		color_arr[2880] = 8'b00010010;
		color_arr[2881] = 8'b00010010;
		color_arr[2882] = 8'b00000000;
		color_arr[2883] = 8'b00000000;
		color_arr[2884] = 8'b00010010;
		color_arr[2885] = 8'b00010010;
		color_arr[2886] = 8'b00010010;
		color_arr[2887] = 8'b00010010;
		color_arr[2888] = 8'b00000010;
		color_arr[2889] = 8'b00000010;
		color_arr[2890] = 8'b00000010;
		color_arr[2891] = 8'b00000010;
		color_arr[2892] = 8'b00000010;
		color_arr[2893] = 8'b00000010;
		color_arr[2894] = 8'b00000010;
		color_arr[2895] = 8'b00000010;
		color_arr[2896] = 8'b00000010;
		color_arr[2897] = 8'b00000010;
		color_arr[2898] = 8'b00000010;
		color_arr[2899] = 8'b00000010;
		color_arr[2900] = 8'b00000010;
		color_arr[2901] = 8'b00000010;
		color_arr[2902] = 8'b00000010;
		color_arr[2903] = 8'b00000010;
		color_arr[2904] = 8'b00000010;
		color_arr[2905] = 8'b00000000;
		color_arr[2906] = 8'b00000000;
		color_arr[2907] = 8'b00000010;
		color_arr[2908] = 8'b00000010;
		color_arr[2909] = 8'b00000010;
		color_arr[2910] = 8'b00000010;
		color_arr[2911] = 8'b00000010;
		color_arr[2912] = 8'b00000010;
		color_arr[2913] = 8'b00000010;
		color_arr[2914] = 8'b00000010;
		color_arr[2915] = 8'b00000010;
		color_arr[2916] = 8'b00000010;
		color_arr[2917] = 8'b00000010;
		color_arr[2918] = 8'b00100000;
		color_arr[2919] = 8'b00100000;
		color_arr[2920] = 8'b00100000;
		color_arr[2921] = 8'b00100000;
		color_arr[2922] = 8'b00100000;
		color_arr[2923] = 8'b00100000;
		color_arr[2924] = 8'b00100000;
		color_arr[2925] = 8'b00100000;
		color_arr[2926] = 8'b00100000;
		color_arr[2927] = 8'b00100000;
		color_arr[2928] = 8'b00100000;
		color_arr[2929] = 8'b00100000;
		color_arr[2930] = 8'b00100000;
		color_arr[2931] = 8'b00100000;
		color_arr[2932] = 8'b00100000;
		color_arr[2933] = 8'b00100000;
		color_arr[2934] = 8'b00100000;
		color_arr[2935] = 8'b00100000;
		color_arr[2936] = 8'b00100000;
		color_arr[2937] = 8'b00100000;
		color_arr[2938] = 8'b00100000;
		color_arr[2939] = 8'b00100000;
		color_arr[2940] = 8'b00100000;
		color_arr[2941] = 8'b00100000;
		color_arr[2942] = 8'b00100000;
		color_arr[2943] = 8'b00100000;
		color_arr[2944] = 8'b00010010;
		color_arr[2945] = 8'b00010010;
		color_arr[2946] = 8'b00000000;
		color_arr[2947] = 8'b00000000;
		color_arr[2948] = 8'b00010010;
		color_arr[2949] = 8'b00010010;
		color_arr[2950] = 8'b00010010;
		color_arr[2951] = 8'b00010010;
		color_arr[2952] = 8'b00000010;
		color_arr[2953] = 8'b00000010;
		color_arr[2954] = 8'b00000010;
		color_arr[2955] = 8'b00000010;
		color_arr[2956] = 8'b00000010;
		color_arr[2957] = 8'b00000010;
		color_arr[2958] = 8'b00000010;
		color_arr[2959] = 8'b00000010;
		color_arr[2960] = 8'b00000010;
		color_arr[2961] = 8'b00000010;
		color_arr[2962] = 8'b00000010;
		color_arr[2963] = 8'b00000010;
		color_arr[2964] = 8'b00000010;
		color_arr[2965] = 8'b00000010;
		color_arr[2966] = 8'b00000010;
		color_arr[2967] = 8'b00000010;
		color_arr[2968] = 8'b00000000;
		color_arr[2969] = 8'b00000000;
		color_arr[2970] = 8'b00000000;
		color_arr[2971] = 8'b00000010;
		color_arr[2972] = 8'b00000010;
		color_arr[2973] = 8'b00000010;
		color_arr[2974] = 8'b00000010;
		color_arr[2975] = 8'b00000010;
		color_arr[2976] = 8'b00000010;
		color_arr[2977] = 8'b00000010;
		color_arr[2978] = 8'b00000010;
		color_arr[2979] = 8'b00000010;
		color_arr[2980] = 8'b00000010;
		color_arr[2981] = 8'b00000010;
		color_arr[2982] = 8'b00100000;
		color_arr[2983] = 8'b00100000;
		color_arr[2984] = 8'b00100000;
		color_arr[2985] = 8'b00100000;
		color_arr[2986] = 8'b00100000;
		color_arr[2987] = 8'b00100000;
		color_arr[2988] = 8'b00100000;
		color_arr[2989] = 8'b00100000;
		color_arr[2990] = 8'b00100000;
		color_arr[2991] = 8'b00100000;
		color_arr[2992] = 8'b00100000;
		color_arr[2993] = 8'b00100000;
		color_arr[2994] = 8'b00100000;
		color_arr[2995] = 8'b00100000;
		color_arr[2996] = 8'b00100000;
		color_arr[2997] = 8'b00100000;
		color_arr[2998] = 8'b00100000;
		color_arr[2999] = 8'b00100000;
		color_arr[3000] = 8'b00100000;
		color_arr[3001] = 8'b00100000;
		color_arr[3002] = 8'b00100000;
		color_arr[3003] = 8'b00100000;
		color_arr[3004] = 8'b00100000;
		color_arr[3005] = 8'b00100000;
		color_arr[3006] = 8'b00100000;
		color_arr[3007] = 8'b00100000;
		color_arr[3008] = 8'b00010010;
		color_arr[3009] = 8'b00010010;
		color_arr[3010] = 8'b00000000;
		color_arr[3011] = 8'b00000000;
		color_arr[3012] = 8'b00010010;
		color_arr[3013] = 8'b00010010;
		color_arr[3014] = 8'b00010010;
		color_arr[3015] = 8'b00010010;
		color_arr[3016] = 8'b00000010;
		color_arr[3017] = 8'b00000010;
		color_arr[3018] = 8'b00000010;
		color_arr[3019] = 8'b00000010;
		color_arr[3020] = 8'b00000010;
		color_arr[3021] = 8'b00000010;
		color_arr[3022] = 8'b00000010;
		color_arr[3023] = 8'b00000010;
		color_arr[3024] = 8'b00000010;
		color_arr[3025] = 8'b00000010;
		color_arr[3026] = 8'b00000010;
		color_arr[3027] = 8'b00000010;
		color_arr[3028] = 8'b00000010;
		color_arr[3029] = 8'b00000010;
		color_arr[3030] = 8'b00000010;
		color_arr[3031] = 8'b00000010;
		color_arr[3032] = 8'b00000000;
		color_arr[3033] = 8'b00000000;
		color_arr[3034] = 8'b00000010;
		color_arr[3035] = 8'b00000010;
		color_arr[3036] = 8'b00000010;
		color_arr[3037] = 8'b00000010;
		color_arr[3038] = 8'b00000010;
		color_arr[3039] = 8'b00000010;
		color_arr[3040] = 8'b00000010;
		color_arr[3041] = 8'b00000010;
		color_arr[3042] = 8'b00000010;
		color_arr[3043] = 8'b00000010;
		color_arr[3044] = 8'b00000010;
		color_arr[3045] = 8'b00000010;
		color_arr[3046] = 8'b00100000;
		color_arr[3047] = 8'b00100000;
		color_arr[3048] = 8'b00100000;
		color_arr[3049] = 8'b00100000;
		color_arr[3050] = 8'b00100000;
		color_arr[3051] = 8'b00100000;
		color_arr[3052] = 8'b00100000;
		color_arr[3053] = 8'b00100000;
		color_arr[3054] = 8'b00100000;
		color_arr[3055] = 8'b00100000;
		color_arr[3056] = 8'b00100000;
		color_arr[3057] = 8'b00100000;
		color_arr[3058] = 8'b00100000;
		color_arr[3059] = 8'b00100000;
		color_arr[3060] = 8'b00100000;
		color_arr[3061] = 8'b00100000;
		color_arr[3062] = 8'b00100000;
		color_arr[3063] = 8'b00100000;
		color_arr[3064] = 8'b00100000;
		color_arr[3065] = 8'b00100000;
		color_arr[3066] = 8'b00100000;
		color_arr[3067] = 8'b00100000;
		color_arr[3068] = 8'b00100000;
		color_arr[3069] = 8'b00100000;
		color_arr[3070] = 8'b00100000;
		color_arr[3071] = 8'b00100000;
		color_arr[3072] = 8'b00010010;
		color_arr[3073] = 8'b00010010;
		color_arr[3074] = 8'b00000000;
		color_arr[3075] = 8'b00000000;
		color_arr[3076] = 8'b00010010;
		color_arr[3077] = 8'b00010010;
		color_arr[3078] = 8'b00010010;
		color_arr[3079] = 8'b00010010;
		color_arr[3080] = 8'b00000010;
		color_arr[3081] = 8'b00000010;
		color_arr[3082] = 8'b00000010;
		color_arr[3083] = 8'b00000010;
		color_arr[3084] = 8'b00000010;
		color_arr[3085] = 8'b00000010;
		color_arr[3086] = 8'b00000010;
		color_arr[3087] = 8'b00000010;
		color_arr[3088] = 8'b00000010;
		color_arr[3089] = 8'b00000010;
		color_arr[3090] = 8'b00000010;
		color_arr[3091] = 8'b00000010;
		color_arr[3092] = 8'b00000010;
		color_arr[3093] = 8'b00000010;
		color_arr[3094] = 8'b00000010;
		color_arr[3095] = 8'b00000000;
		color_arr[3096] = 8'b00000000;
		color_arr[3097] = 8'b00000000;
		color_arr[3098] = 8'b00000010;
		color_arr[3099] = 8'b00000010;
		color_arr[3100] = 8'b00000010;
		color_arr[3101] = 8'b00000010;
		color_arr[3102] = 8'b00000010;
		color_arr[3103] = 8'b00000010;
		color_arr[3104] = 8'b00000010;
		color_arr[3105] = 8'b00000010;
		color_arr[3106] = 8'b00000010;
		color_arr[3107] = 8'b00000010;
		color_arr[3108] = 8'b00000010;
		color_arr[3109] = 8'b00000010;
		color_arr[3110] = 8'b00100000;
		color_arr[3111] = 8'b00100000;
		color_arr[3112] = 8'b00100000;
		color_arr[3113] = 8'b00100000;
		color_arr[3114] = 8'b00100000;
		color_arr[3115] = 8'b00100000;
		color_arr[3116] = 8'b00100000;
		color_arr[3117] = 8'b00100000;
		color_arr[3118] = 8'b00100000;
		color_arr[3119] = 8'b00100000;
		color_arr[3120] = 8'b00100000;
		color_arr[3121] = 8'b00100000;
		color_arr[3122] = 8'b00100000;
		color_arr[3123] = 8'b00100000;
		color_arr[3124] = 8'b00100000;
		color_arr[3125] = 8'b00100000;
		color_arr[3126] = 8'b00100000;
		color_arr[3127] = 8'b00100000;
		color_arr[3128] = 8'b00100000;
		color_arr[3129] = 8'b00100000;
		color_arr[3130] = 8'b00100000;
		color_arr[3131] = 8'b00100000;
		color_arr[3132] = 8'b00100000;
		color_arr[3133] = 8'b00100000;
		color_arr[3134] = 8'b00100000;
		color_arr[3135] = 8'b00100000;
		color_arr[3136] = 8'b00010010;
		color_arr[3137] = 8'b00010010;
		color_arr[3138] = 8'b00000000;
		color_arr[3139] = 8'b00000000;
		color_arr[3140] = 8'b00010010;
		color_arr[3141] = 8'b00010010;
		color_arr[3142] = 8'b00010010;
		color_arr[3143] = 8'b00010010;
		color_arr[3144] = 8'b00000010;
		color_arr[3145] = 8'b00000010;
		color_arr[3146] = 8'b00000010;
		color_arr[3147] = 8'b00000010;
		color_arr[3148] = 8'b00000010;
		color_arr[3149] = 8'b00000010;
		color_arr[3150] = 8'b00000010;
		color_arr[3151] = 8'b00000010;
		color_arr[3152] = 8'b00000010;
		color_arr[3153] = 8'b00000010;
		color_arr[3154] = 8'b00000010;
		color_arr[3155] = 8'b00000010;
		color_arr[3156] = 8'b00000010;
		color_arr[3157] = 8'b00000010;
		color_arr[3158] = 8'b00000010;
		color_arr[3159] = 8'b00000000;
		color_arr[3160] = 8'b00000000;
		color_arr[3161] = 8'b00000010;
		color_arr[3162] = 8'b00000010;
		color_arr[3163] = 8'b00000010;
		color_arr[3164] = 8'b00000010;
		color_arr[3165] = 8'b00000010;
		color_arr[3166] = 8'b00000010;
		color_arr[3167] = 8'b00000010;
		color_arr[3168] = 8'b00000010;
		color_arr[3169] = 8'b00000010;
		color_arr[3170] = 8'b00000010;
		color_arr[3171] = 8'b00000010;
		color_arr[3172] = 8'b00000010;
		color_arr[3173] = 8'b00000010;
		color_arr[3174] = 8'b00100000;
		color_arr[3175] = 8'b00100000;
		color_arr[3176] = 8'b00100000;
		color_arr[3177] = 8'b00100000;
		color_arr[3178] = 8'b00100000;
		color_arr[3179] = 8'b00100000;
		color_arr[3180] = 8'b00100000;
		color_arr[3181] = 8'b00100000;
		color_arr[3182] = 8'b00100000;
		color_arr[3183] = 8'b00100000;
		color_arr[3184] = 8'b00100000;
		color_arr[3185] = 8'b00100000;
		color_arr[3186] = 8'b00100000;
		color_arr[3187] = 8'b00100000;
		color_arr[3188] = 8'b00100000;
		color_arr[3189] = 8'b00100000;
		color_arr[3190] = 8'b00100000;
		color_arr[3191] = 8'b00100000;
		color_arr[3192] = 8'b00100000;
		color_arr[3193] = 8'b00100000;
		color_arr[3194] = 8'b00100000;
		color_arr[3195] = 8'b00100000;
		color_arr[3196] = 8'b00100000;
		color_arr[3197] = 8'b00100000;
		color_arr[3198] = 8'b00100000;
		color_arr[3199] = 8'b00100000;
		color_arr[3200] = 8'b00010010;
		color_arr[3201] = 8'b00010010;
		color_arr[3202] = 8'b00000000;
		color_arr[3203] = 8'b00000000;
		color_arr[3204] = 8'b00010010;
		color_arr[3205] = 8'b00010010;
		color_arr[3206] = 8'b00010010;
		color_arr[3207] = 8'b00010010;
		color_arr[3208] = 8'b00000010;
		color_arr[3209] = 8'b00000010;
		color_arr[3210] = 8'b00000010;
		color_arr[3211] = 8'b00000010;
		color_arr[3212] = 8'b00000010;
		color_arr[3213] = 8'b00000010;
		color_arr[3214] = 8'b00000010;
		color_arr[3215] = 8'b00000010;
		color_arr[3216] = 8'b00000010;
		color_arr[3217] = 8'b00000010;
		color_arr[3218] = 8'b00000010;
		color_arr[3219] = 8'b00000010;
		color_arr[3220] = 8'b00000010;
		color_arr[3221] = 8'b00000010;
		color_arr[3222] = 8'b00000000;
		color_arr[3223] = 8'b00000000;
		color_arr[3224] = 8'b00000000;
		color_arr[3225] = 8'b00000010;
		color_arr[3226] = 8'b00000010;
		color_arr[3227] = 8'b00000010;
		color_arr[3228] = 8'b00000010;
		color_arr[3229] = 8'b00000010;
		color_arr[3230] = 8'b00000010;
		color_arr[3231] = 8'b00000010;
		color_arr[3232] = 8'b00000010;
		color_arr[3233] = 8'b00000010;
		color_arr[3234] = 8'b00000010;
		color_arr[3235] = 8'b00000010;
		color_arr[3236] = 8'b00000010;
		color_arr[3237] = 8'b00000010;
		color_arr[3238] = 8'b00100000;
		color_arr[3239] = 8'b00100000;
		color_arr[3240] = 8'b00100000;
		color_arr[3241] = 8'b00100000;
		color_arr[3242] = 8'b00100000;
		color_arr[3243] = 8'b00100000;
		color_arr[3244] = 8'b00100000;
		color_arr[3245] = 8'b00100000;
		color_arr[3246] = 8'b00100000;
		color_arr[3247] = 8'b00100000;
		color_arr[3248] = 8'b00100000;
		color_arr[3249] = 8'b00100000;
		color_arr[3250] = 8'b00100000;
		color_arr[3251] = 8'b00100000;
		color_arr[3252] = 8'b00100000;
		color_arr[3253] = 8'b00100000;
		color_arr[3254] = 8'b00100000;
		color_arr[3255] = 8'b00100000;
		color_arr[3256] = 8'b00100000;
		color_arr[3257] = 8'b00100000;
		color_arr[3258] = 8'b00100000;
		color_arr[3259] = 8'b00100000;
		color_arr[3260] = 8'b00100000;
		color_arr[3261] = 8'b00100000;
		color_arr[3262] = 8'b00100000;
		color_arr[3263] = 8'b00100000;
		color_arr[3264] = 8'b00010010;
		color_arr[3265] = 8'b00010010;
		color_arr[3266] = 8'b00000000;
		color_arr[3267] = 8'b00000000;
		color_arr[3268] = 8'b00010010;
		color_arr[3269] = 8'b00010010;
		color_arr[3270] = 8'b00010010;
		color_arr[3271] = 8'b00010010;
		color_arr[3272] = 8'b00000010;
		color_arr[3273] = 8'b00000010;
		color_arr[3274] = 8'b00000010;
		color_arr[3275] = 8'b00000010;
		color_arr[3276] = 8'b00000010;
		color_arr[3277] = 8'b00000010;
		color_arr[3278] = 8'b00000010;
		color_arr[3279] = 8'b00000010;
		color_arr[3280] = 8'b00000010;
		color_arr[3281] = 8'b00000010;
		color_arr[3282] = 8'b00000010;
		color_arr[3283] = 8'b00000010;
		color_arr[3284] = 8'b00000010;
		color_arr[3285] = 8'b00000010;
		color_arr[3286] = 8'b00000000;
		color_arr[3287] = 8'b00000000;
		color_arr[3288] = 8'b00000010;
		color_arr[3289] = 8'b00000010;
		color_arr[3290] = 8'b00000010;
		color_arr[3291] = 8'b00000010;
		color_arr[3292] = 8'b00000010;
		color_arr[3293] = 8'b00000010;
		color_arr[3294] = 8'b00000010;
		color_arr[3295] = 8'b00000010;
		color_arr[3296] = 8'b00000010;
		color_arr[3297] = 8'b00000010;
		color_arr[3298] = 8'b00000010;
		color_arr[3299] = 8'b00000010;
		color_arr[3300] = 8'b00000010;
		color_arr[3301] = 8'b00000010;
		color_arr[3302] = 8'b00100000;
		color_arr[3303] = 8'b00100000;
		color_arr[3304] = 8'b00100000;
		color_arr[3305] = 8'b00100000;
		color_arr[3306] = 8'b00100000;
		color_arr[3307] = 8'b00100000;
		color_arr[3308] = 8'b00100000;
		color_arr[3309] = 8'b00100000;
		color_arr[3310] = 8'b00100000;
		color_arr[3311] = 8'b00100000;
		color_arr[3312] = 8'b00100000;
		color_arr[3313] = 8'b00100000;
		color_arr[3314] = 8'b00100000;
		color_arr[3315] = 8'b00100000;
		color_arr[3316] = 8'b00100000;
		color_arr[3317] = 8'b00100000;
		color_arr[3318] = 8'b00100000;
		color_arr[3319] = 8'b00100000;
		color_arr[3320] = 8'b00100000;
		color_arr[3321] = 8'b00100000;
		color_arr[3322] = 8'b00100000;
		color_arr[3323] = 8'b00100000;
		color_arr[3324] = 8'b00100000;
		color_arr[3325] = 8'b00100000;
		color_arr[3326] = 8'b00100000;
		color_arr[3327] = 8'b00100000;
		color_arr[3328] = 8'b00010010;
		color_arr[3329] = 8'b00010010;
		color_arr[3330] = 8'b00000000;
		color_arr[3331] = 8'b00000000;
		color_arr[3332] = 8'b00010010;
		color_arr[3333] = 8'b00010010;
		color_arr[3334] = 8'b00010010;
		color_arr[3335] = 8'b00010010;
		color_arr[3336] = 8'b00000010;
		color_arr[3337] = 8'b00000010;
		color_arr[3338] = 8'b00000010;
		color_arr[3339] = 8'b00000010;
		color_arr[3340] = 8'b00000010;
		color_arr[3341] = 8'b00000010;
		color_arr[3342] = 8'b00000010;
		color_arr[3343] = 8'b00000010;
		color_arr[3344] = 8'b00000010;
		color_arr[3345] = 8'b00000010;
		color_arr[3346] = 8'b00000010;
		color_arr[3347] = 8'b00000010;
		color_arr[3348] = 8'b00000010;
		color_arr[3349] = 8'b00000010;
		color_arr[3350] = 8'b00000000;
		color_arr[3351] = 8'b00000000;
		color_arr[3352] = 8'b00000010;
		color_arr[3353] = 8'b00000010;
		color_arr[3354] = 8'b00000010;
		color_arr[3355] = 8'b00000010;
		color_arr[3356] = 8'b00000010;
		color_arr[3357] = 8'b00000010;
		color_arr[3358] = 8'b00000010;
		color_arr[3359] = 8'b00000010;
		color_arr[3360] = 8'b00000010;
		color_arr[3361] = 8'b00000010;
		color_arr[3362] = 8'b00000010;
		color_arr[3363] = 8'b00000010;
		color_arr[3364] = 8'b00000010;
		color_arr[3365] = 8'b00000010;
		color_arr[3366] = 8'b00100000;
		color_arr[3367] = 8'b00100000;
		color_arr[3368] = 8'b00100000;
		color_arr[3369] = 8'b00100000;
		color_arr[3370] = 8'b00100000;
		color_arr[3371] = 8'b00100000;
		color_arr[3372] = 8'b00100000;
		color_arr[3373] = 8'b00100000;
		color_arr[3374] = 8'b00100000;
		color_arr[3375] = 8'b00100000;
		color_arr[3376] = 8'b00100000;
		color_arr[3377] = 8'b00100000;
		color_arr[3378] = 8'b00100000;
		color_arr[3379] = 8'b00100000;
		color_arr[3380] = 8'b00100000;
		color_arr[3381] = 8'b00100000;
		color_arr[3382] = 8'b00100000;
		color_arr[3383] = 8'b00100000;
		color_arr[3384] = 8'b00100000;
		color_arr[3385] = 8'b00100000;
		color_arr[3386] = 8'b00100000;
		color_arr[3387] = 8'b00100000;
		color_arr[3388] = 8'b00100000;
		color_arr[3389] = 8'b00100000;
		color_arr[3390] = 8'b00100000;
		color_arr[3391] = 8'b00100000;
		color_arr[3392] = 8'b00010010;
		color_arr[3393] = 8'b00010010;
		color_arr[3394] = 8'b00000000;
		color_arr[3395] = 8'b00000000;
		color_arr[3396] = 8'b00010010;
		color_arr[3397] = 8'b00010010;
		color_arr[3398] = 8'b00010010;
		color_arr[3399] = 8'b00010010;
		color_arr[3400] = 8'b00000010;
		color_arr[3401] = 8'b00000010;
		color_arr[3402] = 8'b00000010;
		color_arr[3403] = 8'b00000010;
		color_arr[3404] = 8'b00000010;
		color_arr[3405] = 8'b00000010;
		color_arr[3406] = 8'b00000010;
		color_arr[3407] = 8'b00000010;
		color_arr[3408] = 8'b00000010;
		color_arr[3409] = 8'b00000010;
		color_arr[3410] = 8'b00000010;
		color_arr[3411] = 8'b00000010;
		color_arr[3412] = 8'b00000010;
		color_arr[3413] = 8'b00000010;
		color_arr[3414] = 8'b00000000;
		color_arr[3415] = 8'b00000000;
		color_arr[3416] = 8'b00000010;
		color_arr[3417] = 8'b00000010;
		color_arr[3418] = 8'b00000010;
		color_arr[3419] = 8'b00000010;
		color_arr[3420] = 8'b00000010;
		color_arr[3421] = 8'b00000010;
		color_arr[3422] = 8'b00000010;
		color_arr[3423] = 8'b00000010;
		color_arr[3424] = 8'b00000010;
		color_arr[3425] = 8'b00000010;
		color_arr[3426] = 8'b00000010;
		color_arr[3427] = 8'b00000010;
		color_arr[3428] = 8'b00000010;
		color_arr[3429] = 8'b00000010;
		color_arr[3430] = 8'b00100000;
		color_arr[3431] = 8'b00100000;
		color_arr[3432] = 8'b00100000;
		color_arr[3433] = 8'b00100000;
		color_arr[3434] = 8'b00100000;
		color_arr[3435] = 8'b00100000;
		color_arr[3436] = 8'b00100000;
		color_arr[3437] = 8'b00100000;
		color_arr[3438] = 8'b00100000;
		color_arr[3439] = 8'b00100000;
		color_arr[3440] = 8'b00100000;
		color_arr[3441] = 8'b00100000;
		color_arr[3442] = 8'b00100000;
		color_arr[3443] = 8'b00100000;
		color_arr[3444] = 8'b00100000;
		color_arr[3445] = 8'b00100000;
		color_arr[3446] = 8'b00100000;
		color_arr[3447] = 8'b00100000;
		color_arr[3448] = 8'b00100000;
		color_arr[3449] = 8'b00100000;
		color_arr[3450] = 8'b00100000;
		color_arr[3451] = 8'b00100000;
		color_arr[3452] = 8'b00100000;
		color_arr[3453] = 8'b00100000;
		color_arr[3454] = 8'b00100000;
		color_arr[3455] = 8'b00100000;
		color_arr[3456] = 8'b00010010;
		color_arr[3457] = 8'b00010010;
		color_arr[3458] = 8'b00000000;
		color_arr[3459] = 8'b00000000;
		color_arr[3460] = 8'b00010010;
		color_arr[3461] = 8'b00010010;
		color_arr[3462] = 8'b00010010;
		color_arr[3463] = 8'b00010010;
		color_arr[3464] = 8'b00000010;
		color_arr[3465] = 8'b00000010;
		color_arr[3466] = 8'b00000010;
		color_arr[3467] = 8'b00000010;
		color_arr[3468] = 8'b00000010;
		color_arr[3469] = 8'b00000010;
		color_arr[3470] = 8'b00000010;
		color_arr[3471] = 8'b00000010;
		color_arr[3472] = 8'b00000010;
		color_arr[3473] = 8'b00000010;
		color_arr[3474] = 8'b00000010;
		color_arr[3475] = 8'b00000010;
		color_arr[3476] = 8'b00000010;
		color_arr[3477] = 8'b00000010;
		color_arr[3478] = 8'b00000000;
		color_arr[3479] = 8'b00000000;
		color_arr[3480] = 8'b00000010;
		color_arr[3481] = 8'b00000010;
		color_arr[3482] = 8'b00000010;
		color_arr[3483] = 8'b00000010;
		color_arr[3484] = 8'b00000010;
		color_arr[3485] = 8'b00000010;
		color_arr[3486] = 8'b00000010;
		color_arr[3487] = 8'b00000010;
		color_arr[3488] = 8'b00000010;
		color_arr[3489] = 8'b00000010;
		color_arr[3490] = 8'b00000010;
		color_arr[3491] = 8'b00000010;
		color_arr[3492] = 8'b00000010;
		color_arr[3493] = 8'b00000010;
		color_arr[3494] = 8'b00100000;
		color_arr[3495] = 8'b00100000;
		color_arr[3496] = 8'b00100000;
		color_arr[3497] = 8'b00100000;
		color_arr[3498] = 8'b00100000;
		color_arr[3499] = 8'b00100000;
		color_arr[3500] = 8'b00100000;
		color_arr[3501] = 8'b00100000;
		color_arr[3502] = 8'b00100000;
		color_arr[3503] = 8'b00100000;
		color_arr[3504] = 8'b00100000;
		color_arr[3505] = 8'b00100000;
		color_arr[3506] = 8'b00100000;
		color_arr[3507] = 8'b00100000;
		color_arr[3508] = 8'b00100000;
		color_arr[3509] = 8'b00100000;
		color_arr[3510] = 8'b00100000;
		color_arr[3511] = 8'b00100000;
		color_arr[3512] = 8'b00100000;
		color_arr[3513] = 8'b00100000;
		color_arr[3514] = 8'b00100000;
		color_arr[3515] = 8'b00100000;
		color_arr[3516] = 8'b00100000;
		color_arr[3517] = 8'b00100000;
		color_arr[3518] = 8'b00100000;
		color_arr[3519] = 8'b00100000;
		color_arr[3520] = 8'b00010010;
		color_arr[3521] = 8'b00010010;
		color_arr[3522] = 8'b00000000;
		color_arr[3523] = 8'b00000000;
		color_arr[3524] = 8'b00010010;
		color_arr[3525] = 8'b00010010;
		color_arr[3526] = 8'b00010010;
		color_arr[3527] = 8'b00010010;
		color_arr[3528] = 8'b00010010;
		color_arr[3529] = 8'b00010010;
		color_arr[3530] = 8'b00010010;
		color_arr[3531] = 8'b00010010;
		color_arr[3532] = 8'b00010010;
		color_arr[3533] = 8'b00010010;
		color_arr[3534] = 8'b00010010;
		color_arr[3535] = 8'b00010010;
		color_arr[3536] = 8'b00010010;
		color_arr[3537] = 8'b00010010;
		color_arr[3538] = 8'b00100000;
		color_arr[3539] = 8'b00100000;
		color_arr[3540] = 8'b00100000;
		color_arr[3541] = 8'b00100000;
		color_arr[3542] = 8'b00000000;
		color_arr[3543] = 8'b00000000;
		color_arr[3544] = 8'b00100000;
		color_arr[3545] = 8'b00100000;
		color_arr[3546] = 8'b00100000;
		color_arr[3547] = 8'b00100000;
		color_arr[3548] = 8'b00100000;
		color_arr[3549] = 8'b00100000;
		color_arr[3550] = 8'b00100000;
		color_arr[3551] = 8'b00100000;
		color_arr[3552] = 8'b00100000;
		color_arr[3553] = 8'b00100000;
		color_arr[3554] = 8'b00100000;
		color_arr[3555] = 8'b00100000;
		color_arr[3556] = 8'b00100000;
		color_arr[3557] = 8'b00100000;
		color_arr[3558] = 8'b00100000;
		color_arr[3559] = 8'b00100000;
		color_arr[3560] = 8'b00100000;
		color_arr[3561] = 8'b00100000;
		color_arr[3562] = 8'b00100000;
		color_arr[3563] = 8'b00100000;
		color_arr[3564] = 8'b00100000;
		color_arr[3565] = 8'b00100000;
		color_arr[3566] = 8'b00100000;
		color_arr[3567] = 8'b00100000;
		color_arr[3568] = 8'b00100000;
		color_arr[3569] = 8'b00100000;
		color_arr[3570] = 8'b00100000;
		color_arr[3571] = 8'b00100000;
		color_arr[3572] = 8'b00100000;
		color_arr[3573] = 8'b00100000;
		color_arr[3574] = 8'b00100000;
		color_arr[3575] = 8'b00100000;
		color_arr[3576] = 8'b00100000;
		color_arr[3577] = 8'b00100000;
		color_arr[3578] = 8'b00100000;
		color_arr[3579] = 8'b00100000;
		color_arr[3580] = 8'b00100000;
		color_arr[3581] = 8'b00100000;
		color_arr[3582] = 8'b00100000;
		color_arr[3583] = 8'b00100000;
		color_arr[3584] = 8'b00010010;
		color_arr[3585] = 8'b00010010;
		color_arr[3586] = 8'b00000000;
		color_arr[3587] = 8'b00000000;
		color_arr[3588] = 8'b00010010;
		color_arr[3589] = 8'b00010010;
		color_arr[3590] = 8'b00010010;
		color_arr[3591] = 8'b00010010;
		color_arr[3592] = 8'b00010010;
		color_arr[3593] = 8'b00010010;
		color_arr[3594] = 8'b00010010;
		color_arr[3595] = 8'b00010010;
		color_arr[3596] = 8'b00010010;
		color_arr[3597] = 8'b00010010;
		color_arr[3598] = 8'b00010010;
		color_arr[3599] = 8'b00010010;
		color_arr[3600] = 8'b00010010;
		color_arr[3601] = 8'b00010010;
		color_arr[3602] = 8'b00100000;
		color_arr[3603] = 8'b00100000;
		color_arr[3604] = 8'b00100000;
		color_arr[3605] = 8'b00000000;
		color_arr[3606] = 8'b00000000;
		color_arr[3607] = 8'b00000000;
		color_arr[3608] = 8'b00100000;
		color_arr[3609] = 8'b00100000;
		color_arr[3610] = 8'b00100000;
		color_arr[3611] = 8'b00100000;
		color_arr[3612] = 8'b00100000;
		color_arr[3613] = 8'b00100000;
		color_arr[3614] = 8'b00100000;
		color_arr[3615] = 8'b00100000;
		color_arr[3616] = 8'b00100000;
		color_arr[3617] = 8'b00100000;
		color_arr[3618] = 8'b00100000;
		color_arr[3619] = 8'b00100000;
		color_arr[3620] = 8'b00100000;
		color_arr[3621] = 8'b00100000;
		color_arr[3622] = 8'b00100000;
		color_arr[3623] = 8'b00100000;
		color_arr[3624] = 8'b00100000;
		color_arr[3625] = 8'b00100000;
		color_arr[3626] = 8'b00100000;
		color_arr[3627] = 8'b00100000;
		color_arr[3628] = 8'b00100000;
		color_arr[3629] = 8'b00100000;
		color_arr[3630] = 8'b00100000;
		color_arr[3631] = 8'b00100000;
		color_arr[3632] = 8'b00100000;
		color_arr[3633] = 8'b00100000;
		color_arr[3634] = 8'b00100000;
		color_arr[3635] = 8'b00100000;
		color_arr[3636] = 8'b00100000;
		color_arr[3637] = 8'b00100000;
		color_arr[3638] = 8'b00100000;
		color_arr[3639] = 8'b00100000;
		color_arr[3640] = 8'b00100000;
		color_arr[3641] = 8'b00100000;
		color_arr[3642] = 8'b00100000;
		color_arr[3643] = 8'b00100000;
		color_arr[3644] = 8'b00100000;
		color_arr[3645] = 8'b00100000;
		color_arr[3646] = 8'b00100000;
		color_arr[3647] = 8'b00100000;
		color_arr[3648] = 8'b00010010;
		color_arr[3649] = 8'b00010010;
		color_arr[3650] = 8'b00000000;
		color_arr[3651] = 8'b00000000;
		color_arr[3652] = 8'b00010010;
		color_arr[3653] = 8'b00010010;
		color_arr[3654] = 8'b00010010;
		color_arr[3655] = 8'b00010010;
		color_arr[3656] = 8'b00010010;
		color_arr[3657] = 8'b00010010;
		color_arr[3658] = 8'b00010010;
		color_arr[3659] = 8'b00010010;
		color_arr[3660] = 8'b00010010;
		color_arr[3661] = 8'b00010010;
		color_arr[3662] = 8'b00010010;
		color_arr[3663] = 8'b00010010;
		color_arr[3664] = 8'b00010010;
		color_arr[3665] = 8'b00010010;
		color_arr[3666] = 8'b00100000;
		color_arr[3667] = 8'b00100000;
		color_arr[3668] = 8'b00100000;
		color_arr[3669] = 8'b00000000;
		color_arr[3670] = 8'b00000000;
		color_arr[3671] = 8'b00100000;
		color_arr[3672] = 8'b00100000;
		color_arr[3673] = 8'b00100000;
		color_arr[3674] = 8'b00100000;
		color_arr[3675] = 8'b00100000;
		color_arr[3676] = 8'b00100000;
		color_arr[3677] = 8'b00100000;
		color_arr[3678] = 8'b00100000;
		color_arr[3679] = 8'b00100000;
		color_arr[3680] = 8'b00100000;
		color_arr[3681] = 8'b00100000;
		color_arr[3682] = 8'b00100000;
		color_arr[3683] = 8'b00100000;
		color_arr[3684] = 8'b00100000;
		color_arr[3685] = 8'b00100000;
		color_arr[3686] = 8'b00100000;
		color_arr[3687] = 8'b00100000;
		color_arr[3688] = 8'b00100000;
		color_arr[3689] = 8'b00100000;
		color_arr[3690] = 8'b00100000;
		color_arr[3691] = 8'b00100000;
		color_arr[3692] = 8'b00100000;
		color_arr[3693] = 8'b00100000;
		color_arr[3694] = 8'b00100000;
		color_arr[3695] = 8'b00100000;
		color_arr[3696] = 8'b00100000;
		color_arr[3697] = 8'b00100000;
		color_arr[3698] = 8'b00100000;
		color_arr[3699] = 8'b00100000;
		color_arr[3700] = 8'b00100000;
		color_arr[3701] = 8'b00100000;
		color_arr[3702] = 8'b00100000;
		color_arr[3703] = 8'b00100000;
		color_arr[3704] = 8'b00100000;
		color_arr[3705] = 8'b00100000;
		color_arr[3706] = 8'b00100000;
		color_arr[3707] = 8'b00100000;
		color_arr[3708] = 8'b00100000;
		color_arr[3709] = 8'b00100000;
		color_arr[3710] = 8'b00100000;
		color_arr[3711] = 8'b00100000;
		color_arr[3712] = 8'b00010010;
		color_arr[3713] = 8'b00010010;
		color_arr[3714] = 8'b00000000;
		color_arr[3715] = 8'b00000000;
		color_arr[3716] = 8'b00010010;
		color_arr[3717] = 8'b00010010;
		color_arr[3718] = 8'b00010010;
		color_arr[3719] = 8'b00010010;
		color_arr[3720] = 8'b00010010;
		color_arr[3721] = 8'b00010010;
		color_arr[3722] = 8'b00010010;
		color_arr[3723] = 8'b00010010;
		color_arr[3724] = 8'b00010010;
		color_arr[3725] = 8'b00010010;
		color_arr[3726] = 8'b00010010;
		color_arr[3727] = 8'b00010010;
		color_arr[3728] = 8'b00010010;
		color_arr[3729] = 8'b00010010;
		color_arr[3730] = 8'b00100000;
		color_arr[3731] = 8'b00100000;
		color_arr[3732] = 8'b00100000;
		color_arr[3733] = 8'b00000000;
		color_arr[3734] = 8'b00000000;
		color_arr[3735] = 8'b00100000;
		color_arr[3736] = 8'b00100000;
		color_arr[3737] = 8'b00100000;
		color_arr[3738] = 8'b00100000;
		color_arr[3739] = 8'b00100000;
		color_arr[3740] = 8'b00100000;
		color_arr[3741] = 8'b00100000;
		color_arr[3742] = 8'b00100000;
		color_arr[3743] = 8'b00100000;
		color_arr[3744] = 8'b00100000;
		color_arr[3745] = 8'b00100000;
		color_arr[3746] = 8'b00100000;
		color_arr[3747] = 8'b00100000;
		color_arr[3748] = 8'b00100000;
		color_arr[3749] = 8'b00100000;
		color_arr[3750] = 8'b00100000;
		color_arr[3751] = 8'b00100000;
		color_arr[3752] = 8'b00100000;
		color_arr[3753] = 8'b00100000;
		color_arr[3754] = 8'b00100000;
		color_arr[3755] = 8'b00100000;
		color_arr[3756] = 8'b00100000;
		color_arr[3757] = 8'b00100000;
		color_arr[3758] = 8'b00100000;
		color_arr[3759] = 8'b00100000;
		color_arr[3760] = 8'b00100000;
		color_arr[3761] = 8'b00100000;
		color_arr[3762] = 8'b00100000;
		color_arr[3763] = 8'b00100000;
		color_arr[3764] = 8'b00100000;
		color_arr[3765] = 8'b00100000;
		color_arr[3766] = 8'b00100000;
		color_arr[3767] = 8'b00100000;
		color_arr[3768] = 8'b00100000;
		color_arr[3769] = 8'b00100000;
		color_arr[3770] = 8'b00100000;
		color_arr[3771] = 8'b00100000;
		color_arr[3772] = 8'b00100000;
		color_arr[3773] = 8'b00100000;
		color_arr[3774] = 8'b00100000;
		color_arr[3775] = 8'b00100000;
		color_arr[3776] = 8'b00010010;
		color_arr[3777] = 8'b00010010;
		color_arr[3778] = 8'b00000000;
		color_arr[3779] = 8'b00000000;
		color_arr[3780] = 8'b00010010;
		color_arr[3781] = 8'b00010010;
		color_arr[3782] = 8'b00010010;
		color_arr[3783] = 8'b00010010;
		color_arr[3784] = 8'b00010010;
		color_arr[3785] = 8'b00010010;
		color_arr[3786] = 8'b00010010;
		color_arr[3787] = 8'b00010010;
		color_arr[3788] = 8'b00010010;
		color_arr[3789] = 8'b00010010;
		color_arr[3790] = 8'b00010010;
		color_arr[3791] = 8'b00010010;
		color_arr[3792] = 8'b00010010;
		color_arr[3793] = 8'b00010010;
		color_arr[3794] = 8'b00100000;
		color_arr[3795] = 8'b00100000;
		color_arr[3796] = 8'b00100000;
		color_arr[3797] = 8'b00000000;
		color_arr[3798] = 8'b00000000;
		color_arr[3799] = 8'b00100000;
		color_arr[3800] = 8'b00100000;
		color_arr[3801] = 8'b00100000;
		color_arr[3802] = 8'b00100000;
		color_arr[3803] = 8'b00100000;
		color_arr[3804] = 8'b00100000;
		color_arr[3805] = 8'b00100000;
		color_arr[3806] = 8'b00100000;
		color_arr[3807] = 8'b00100000;
		color_arr[3808] = 8'b00100000;
		color_arr[3809] = 8'b00100000;
		color_arr[3810] = 8'b00100000;
		color_arr[3811] = 8'b00100000;
		color_arr[3812] = 8'b00100000;
		color_arr[3813] = 8'b00100000;
		color_arr[3814] = 8'b00100000;
		color_arr[3815] = 8'b00100000;
		color_arr[3816] = 8'b00100000;
		color_arr[3817] = 8'b00100000;
		color_arr[3818] = 8'b00100000;
		color_arr[3819] = 8'b00100000;
		color_arr[3820] = 8'b00100000;
		color_arr[3821] = 8'b00100000;
		color_arr[3822] = 8'b00100000;
		color_arr[3823] = 8'b00100000;
		color_arr[3824] = 8'b00100000;
		color_arr[3825] = 8'b00100000;
		color_arr[3826] = 8'b00100000;
		color_arr[3827] = 8'b00100000;
		color_arr[3828] = 8'b00100000;
		color_arr[3829] = 8'b00100000;
		color_arr[3830] = 8'b00100000;
		color_arr[3831] = 8'b00100000;
		color_arr[3832] = 8'b00100000;
		color_arr[3833] = 8'b00100000;
		color_arr[3834] = 8'b00100000;
		color_arr[3835] = 8'b00100000;
		color_arr[3836] = 8'b00100000;
		color_arr[3837] = 8'b00100000;
		color_arr[3838] = 8'b00100000;
		color_arr[3839] = 8'b00100000;
		color_arr[3840] = 8'b00010010;
		color_arr[3841] = 8'b00010010;
		color_arr[3842] = 8'b00000000;
		color_arr[3843] = 8'b00000000;
		color_arr[3844] = 8'b00010010;
		color_arr[3845] = 8'b00010010;
		color_arr[3846] = 8'b00010010;
		color_arr[3847] = 8'b00010010;
		color_arr[3848] = 8'b00010010;
		color_arr[3849] = 8'b00010010;
		color_arr[3850] = 8'b00010010;
		color_arr[3851] = 8'b00010010;
		color_arr[3852] = 8'b00010010;
		color_arr[3853] = 8'b00010010;
		color_arr[3854] = 8'b00010010;
		color_arr[3855] = 8'b00010010;
		color_arr[3856] = 8'b00010010;
		color_arr[3857] = 8'b00010010;
		color_arr[3858] = 8'b00100000;
		color_arr[3859] = 8'b00100000;
		color_arr[3860] = 8'b00100000;
		color_arr[3861] = 8'b00000000;
		color_arr[3862] = 8'b00000000;
		color_arr[3863] = 8'b00100000;
		color_arr[3864] = 8'b00100000;
		color_arr[3865] = 8'b00100000;
		color_arr[3866] = 8'b00100000;
		color_arr[3867] = 8'b00100000;
		color_arr[3868] = 8'b00100000;
		color_arr[3869] = 8'b00100000;
		color_arr[3870] = 8'b00100000;
		color_arr[3871] = 8'b00100000;
		color_arr[3872] = 8'b00100000;
		color_arr[3873] = 8'b00100000;
		color_arr[3874] = 8'b00100000;
		color_arr[3875] = 8'b00100000;
		color_arr[3876] = 8'b00100000;
		color_arr[3877] = 8'b00100000;
		color_arr[3878] = 8'b00100000;
		color_arr[3879] = 8'b00100000;
		color_arr[3880] = 8'b00100000;
		color_arr[3881] = 8'b00100000;
		color_arr[3882] = 8'b00100000;
		color_arr[3883] = 8'b00100000;
		color_arr[3884] = 8'b00100000;
		color_arr[3885] = 8'b00100000;
		color_arr[3886] = 8'b00100000;
		color_arr[3887] = 8'b00100000;
		color_arr[3888] = 8'b00100000;
		color_arr[3889] = 8'b00100000;
		color_arr[3890] = 8'b00100000;
		color_arr[3891] = 8'b00100000;
		color_arr[3892] = 8'b00100000;
		color_arr[3893] = 8'b00100000;
		color_arr[3894] = 8'b00100000;
		color_arr[3895] = 8'b00100000;
		color_arr[3896] = 8'b00100000;
		color_arr[3897] = 8'b00100000;
		color_arr[3898] = 8'b00100000;
		color_arr[3899] = 8'b00100000;
		color_arr[3900] = 8'b00100000;
		color_arr[3901] = 8'b00100000;
		color_arr[3902] = 8'b00100000;
		color_arr[3903] = 8'b00100000;
		color_arr[3904] = 8'b00010010;
		color_arr[3905] = 8'b00010010;
		color_arr[3906] = 8'b00000000;
		color_arr[3907] = 8'b00000000;
		color_arr[3908] = 8'b00010010;
		color_arr[3909] = 8'b00010010;
		color_arr[3910] = 8'b00010010;
		color_arr[3911] = 8'b00010010;
		color_arr[3912] = 8'b00010010;
		color_arr[3913] = 8'b00010010;
		color_arr[3914] = 8'b00010010;
		color_arr[3915] = 8'b00010010;
		color_arr[3916] = 8'b00010010;
		color_arr[3917] = 8'b00010010;
		color_arr[3918] = 8'b00010010;
		color_arr[3919] = 8'b00010010;
		color_arr[3920] = 8'b00010010;
		color_arr[3921] = 8'b00010010;
		color_arr[3922] = 8'b00100000;
		color_arr[3923] = 8'b00100000;
		color_arr[3924] = 8'b00100000;
		color_arr[3925] = 8'b00000000;
		color_arr[3926] = 8'b00000000;
		color_arr[3927] = 8'b00100000;
		color_arr[3928] = 8'b00100000;
		color_arr[3929] = 8'b00100000;
		color_arr[3930] = 8'b00100000;
		color_arr[3931] = 8'b00100000;
		color_arr[3932] = 8'b00100000;
		color_arr[3933] = 8'b00100000;
		color_arr[3934] = 8'b00100000;
		color_arr[3935] = 8'b00100000;
		color_arr[3936] = 8'b00100000;
		color_arr[3937] = 8'b00100000;
		color_arr[3938] = 8'b00100000;
		color_arr[3939] = 8'b00100000;
		color_arr[3940] = 8'b00100000;
		color_arr[3941] = 8'b00100000;
		color_arr[3942] = 8'b00100000;
		color_arr[3943] = 8'b00100000;
		color_arr[3944] = 8'b00100000;
		color_arr[3945] = 8'b00100000;
		color_arr[3946] = 8'b00100000;
		color_arr[3947] = 8'b00100000;
		color_arr[3948] = 8'b00100000;
		color_arr[3949] = 8'b00100000;
		color_arr[3950] = 8'b00100000;
		color_arr[3951] = 8'b00100000;
		color_arr[3952] = 8'b00100000;
		color_arr[3953] = 8'b00100000;
		color_arr[3954] = 8'b00100000;
		color_arr[3955] = 8'b00100000;
		color_arr[3956] = 8'b00100000;
		color_arr[3957] = 8'b00100000;
		color_arr[3958] = 8'b00100000;
		color_arr[3959] = 8'b00100000;
		color_arr[3960] = 8'b00100000;
		color_arr[3961] = 8'b00100000;
		color_arr[3962] = 8'b00100000;
		color_arr[3963] = 8'b00100000;
		color_arr[3964] = 8'b00100000;
		color_arr[3965] = 8'b00100000;
		color_arr[3966] = 8'b00100000;
		color_arr[3967] = 8'b00100000;
		color_arr[3968] = 8'b00010010;
		color_arr[3969] = 8'b00010010;
		color_arr[3970] = 8'b00000000;
		color_arr[3971] = 8'b00000000;
		color_arr[3972] = 8'b00010010;
		color_arr[3973] = 8'b00010010;
		color_arr[3974] = 8'b00010010;
		color_arr[3975] = 8'b00010010;
		color_arr[3976] = 8'b00010010;
		color_arr[3977] = 8'b00010010;
		color_arr[3978] = 8'b00010010;
		color_arr[3979] = 8'b00010010;
		color_arr[3980] = 8'b00010010;
		color_arr[3981] = 8'b00010010;
		color_arr[3982] = 8'b00010010;
		color_arr[3983] = 8'b00010010;
		color_arr[3984] = 8'b00010010;
		color_arr[3985] = 8'b00010010;
		color_arr[3986] = 8'b00100000;
		color_arr[3987] = 8'b00100000;
		color_arr[3988] = 8'b00100000;
		color_arr[3989] = 8'b00000000;
		color_arr[3990] = 8'b00000000;
		color_arr[3991] = 8'b00100000;
		color_arr[3992] = 8'b00100000;
		color_arr[3993] = 8'b00100000;
		color_arr[3994] = 8'b00100000;
		color_arr[3995] = 8'b00100000;
		color_arr[3996] = 8'b00100000;
		color_arr[3997] = 8'b00100000;
		color_arr[3998] = 8'b00100000;
		color_arr[3999] = 8'b00100000;
		color_arr[4000] = 8'b00100000;
		color_arr[4001] = 8'b00100000;
		color_arr[4002] = 8'b00100000;
		color_arr[4003] = 8'b00100000;
		color_arr[4004] = 8'b00100000;
		color_arr[4005] = 8'b00100000;
		color_arr[4006] = 8'b00100000;
		color_arr[4007] = 8'b00100000;
		color_arr[4008] = 8'b00100000;
		color_arr[4009] = 8'b00100000;
		color_arr[4010] = 8'b00100000;
		color_arr[4011] = 8'b00100000;
		color_arr[4012] = 8'b00100000;
		color_arr[4013] = 8'b00100000;
		color_arr[4014] = 8'b00100000;
		color_arr[4015] = 8'b00100000;
		color_arr[4016] = 8'b00100000;
		color_arr[4017] = 8'b00100000;
		color_arr[4018] = 8'b00100000;
		color_arr[4019] = 8'b00100000;
		color_arr[4020] = 8'b00100000;
		color_arr[4021] = 8'b00100000;
		color_arr[4022] = 8'b00100000;
		color_arr[4023] = 8'b00100000;
		color_arr[4024] = 8'b00100000;
		color_arr[4025] = 8'b00100000;
		color_arr[4026] = 8'b00100000;
		color_arr[4027] = 8'b00100000;
		color_arr[4028] = 8'b00100000;
		color_arr[4029] = 8'b00100000;
		color_arr[4030] = 8'b00100000;
		color_arr[4031] = 8'b00100000;
		color_arr[4032] = 8'b00010010;
		color_arr[4033] = 8'b00010010;
		color_arr[4034] = 8'b00000000;
		color_arr[4035] = 8'b00000000;
		color_arr[4036] = 8'b00010010;
		color_arr[4037] = 8'b00010010;
		color_arr[4038] = 8'b00010010;
		color_arr[4039] = 8'b00010010;
		color_arr[4040] = 8'b00010010;
		color_arr[4041] = 8'b00010010;
		color_arr[4042] = 8'b00010010;
		color_arr[4043] = 8'b00010010;
		color_arr[4044] = 8'b00010010;
		color_arr[4045] = 8'b00010010;
		color_arr[4046] = 8'b00010010;
		color_arr[4047] = 8'b00010010;
		color_arr[4048] = 8'b00010010;
		color_arr[4049] = 8'b00010010;
		color_arr[4050] = 8'b00100000;
		color_arr[4051] = 8'b00100000;
		color_arr[4052] = 8'b00100000;
		color_arr[4053] = 8'b00000000;
		color_arr[4054] = 8'b00000000;
		color_arr[4055] = 8'b00100000;
		color_arr[4056] = 8'b00100000;
		color_arr[4057] = 8'b00100000;
		color_arr[4058] = 8'b00100000;
		color_arr[4059] = 8'b00100000;
		color_arr[4060] = 8'b00100000;
		color_arr[4061] = 8'b00100000;
		color_arr[4062] = 8'b00100000;
		color_arr[4063] = 8'b00100000;
		color_arr[4064] = 8'b00100000;
		color_arr[4065] = 8'b00100000;
		color_arr[4066] = 8'b00100000;
		color_arr[4067] = 8'b00100000;
		color_arr[4068] = 8'b00100000;
		color_arr[4069] = 8'b00100000;
		color_arr[4070] = 8'b00100000;
		color_arr[4071] = 8'b00100000;
		color_arr[4072] = 8'b00100000;
		color_arr[4073] = 8'b00100000;
		color_arr[4074] = 8'b00100000;
		color_arr[4075] = 8'b00100000;
		color_arr[4076] = 8'b00100000;
		color_arr[4077] = 8'b00100000;
		color_arr[4078] = 8'b00100000;
		color_arr[4079] = 8'b00100000;
		color_arr[4080] = 8'b00100000;
		color_arr[4081] = 8'b00100000;
		color_arr[4082] = 8'b00100000;
		color_arr[4083] = 8'b00100000;
		color_arr[4084] = 8'b00100000;
		color_arr[4085] = 8'b00100000;
		color_arr[4086] = 8'b00100000;
		color_arr[4087] = 8'b00100000;
		color_arr[4088] = 8'b00100000;
		color_arr[4089] = 8'b00100000;
		color_arr[4090] = 8'b00100000;
		color_arr[4091] = 8'b00100000;
		color_arr[4092] = 8'b00100000;
		color_arr[4093] = 8'b00100000;
		color_arr[4094] = 8'b00100000;
		color_arr[4095] = 8'b00100000;
	end

	always @(posedge clk) begin
		color_out <= color_arr[addr][5:0];
	end
endmodule
