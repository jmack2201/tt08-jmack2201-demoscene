module sprite_rom (
	input clk,
	input [13:0] addr,
	output reg [5:0] color_out
);
	reg [7:0] color_arr [SPRITE_SIZE*SPRITE_SIZE-1:0];

	initial begin
		color_arr[0] = 8'b00010010;
		color_arr[1] = 8'b00010010;
		color_arr[2] = 8'b00010010;
		color_arr[3] = 8'b00010010;
		color_arr[4] = 8'b00010010;
		color_arr[5] = 8'b00010010;
		color_arr[6] = 8'b00010010;
		color_arr[7] = 8'b00010010;
		color_arr[8] = 8'b00010010;
		color_arr[9] = 8'b00010010;
		color_arr[10] = 8'b00010010;
		color_arr[11] = 8'b00010010;
		color_arr[12] = 8'b00010010;
		color_arr[13] = 8'b00010010;
		color_arr[14] = 8'b00010010;
		color_arr[15] = 8'b00010010;
		color_arr[16] = 8'b00010010;
		color_arr[17] = 8'b00010010;
		color_arr[18] = 8'b00010010;
		color_arr[19] = 8'b00010010;
		color_arr[20] = 8'b00010010;
		color_arr[21] = 8'b00010010;
		color_arr[22] = 8'b00010010;
		color_arr[23] = 8'b00010010;
		color_arr[24] = 8'b00010010;
		color_arr[25] = 8'b00010010;
		color_arr[26] = 8'b00010010;
		color_arr[27] = 8'b00010010;
		color_arr[28] = 8'b00010010;
		color_arr[29] = 8'b00010010;
		color_arr[30] = 8'b00010010;
		color_arr[31] = 8'b00010010;
		color_arr[32] = 8'b00010010;
		color_arr[33] = 8'b00010010;
		color_arr[34] = 8'b00010010;
		color_arr[35] = 8'b00010010;
		color_arr[36] = 8'b00010010;
		color_arr[37] = 8'b00010010;
		color_arr[38] = 8'b00010010;
		color_arr[39] = 8'b00010010;
		color_arr[40] = 8'b00010010;
		color_arr[41] = 8'b00010010;
		color_arr[42] = 8'b00010010;
		color_arr[43] = 8'b00010010;
		color_arr[44] = 8'b00010010;
		color_arr[45] = 8'b00010010;
		color_arr[46] = 8'b00010010;
		color_arr[47] = 8'b00010010;
		color_arr[48] = 8'b00010010;
		color_arr[49] = 8'b00010010;
		color_arr[50] = 8'b00010010;
		color_arr[51] = 8'b00010010;
		color_arr[52] = 8'b00010010;
		color_arr[53] = 8'b00010010;
		color_arr[54] = 8'b00010010;
		color_arr[55] = 8'b00010010;
		color_arr[56] = 8'b00010010;
		color_arr[57] = 8'b00010010;
		color_arr[58] = 8'b00010010;
		color_arr[59] = 8'b00010010;
		color_arr[60] = 8'b00010010;
		color_arr[61] = 8'b00010010;
		color_arr[62] = 8'b00010010;
		color_arr[63] = 8'b00010010;
		color_arr[64] = 8'b00000000;
		color_arr[65] = 8'b00000000;
		color_arr[66] = 8'b00000000;
		color_arr[67] = 8'b00000000;
		color_arr[68] = 8'b00000000;
		color_arr[69] = 8'b00000000;
		color_arr[70] = 8'b00000000;
		color_arr[71] = 8'b00000000;
		color_arr[72] = 8'b00000000;
		color_arr[73] = 8'b00000000;
		color_arr[74] = 8'b00000000;
		color_arr[75] = 8'b00000000;
		color_arr[76] = 8'b00000000;
		color_arr[77] = 8'b00000000;
		color_arr[78] = 8'b00000000;
		color_arr[79] = 8'b00000000;
		color_arr[80] = 8'b00000000;
		color_arr[81] = 8'b00010010;
		color_arr[82] = 8'b00010010;
		color_arr[83] = 8'b00010010;
		color_arr[84] = 8'b00010010;
		color_arr[85] = 8'b00010010;
		color_arr[86] = 8'b00010010;
		color_arr[87] = 8'b00010010;
		color_arr[88] = 8'b00010010;
		color_arr[89] = 8'b00010010;
		color_arr[90] = 8'b00010010;
		color_arr[91] = 8'b00010010;
		color_arr[92] = 8'b00010010;
		color_arr[93] = 8'b00010010;
		color_arr[94] = 8'b00010010;
		color_arr[95] = 8'b00010010;
		color_arr[96] = 8'b00010010;
		color_arr[97] = 8'b00010010;
		color_arr[98] = 8'b00010010;
		color_arr[99] = 8'b00010010;
		color_arr[100] = 8'b00010010;
		color_arr[101] = 8'b00010010;
		color_arr[102] = 8'b00010010;
		color_arr[103] = 8'b00010010;
		color_arr[104] = 8'b00010010;
		color_arr[105] = 8'b00010010;
		color_arr[106] = 8'b00010010;
		color_arr[107] = 8'b00010010;
		color_arr[108] = 8'b00010010;
		color_arr[109] = 8'b00010010;
		color_arr[110] = 8'b00010010;
		color_arr[111] = 8'b00010010;
		color_arr[112] = 8'b00010010;
		color_arr[113] = 8'b00010010;
		color_arr[114] = 8'b00010010;
		color_arr[115] = 8'b00010010;
		color_arr[116] = 8'b00010010;
		color_arr[117] = 8'b00010010;
		color_arr[118] = 8'b00010010;
		color_arr[119] = 8'b00010010;
		color_arr[120] = 8'b00010010;
		color_arr[121] = 8'b00010010;
		color_arr[122] = 8'b00010010;
		color_arr[123] = 8'b00010010;
		color_arr[124] = 8'b00010010;
		color_arr[125] = 8'b00010010;
		color_arr[126] = 8'b00010010;
		color_arr[127] = 8'b00010010;
		color_arr[128] = 8'b00010010;
		color_arr[129] = 8'b00010010;
		color_arr[130] = 8'b00010010;
		color_arr[131] = 8'b00010010;
		color_arr[132] = 8'b00010010;
		color_arr[133] = 8'b00010010;
		color_arr[134] = 8'b00010010;
		color_arr[135] = 8'b00010010;
		color_arr[136] = 8'b00010010;
		color_arr[137] = 8'b00010010;
		color_arr[138] = 8'b00010010;
		color_arr[139] = 8'b00010010;
		color_arr[140] = 8'b00010010;
		color_arr[141] = 8'b00010010;
		color_arr[142] = 8'b00010010;
		color_arr[143] = 8'b00010010;
		color_arr[144] = 8'b00010010;
		color_arr[145] = 8'b00010010;
		color_arr[146] = 8'b00010010;
		color_arr[147] = 8'b00010010;
		color_arr[148] = 8'b00010010;
		color_arr[149] = 8'b00010010;
		color_arr[150] = 8'b00010010;
		color_arr[151] = 8'b00010010;
		color_arr[152] = 8'b00010010;
		color_arr[153] = 8'b00010010;
		color_arr[154] = 8'b00010010;
		color_arr[155] = 8'b00010010;
		color_arr[156] = 8'b00010010;
		color_arr[157] = 8'b00010010;
		color_arr[158] = 8'b00010010;
		color_arr[159] = 8'b00010010;
		color_arr[160] = 8'b00010010;
		color_arr[161] = 8'b00010010;
		color_arr[162] = 8'b00010010;
		color_arr[163] = 8'b00010010;
		color_arr[164] = 8'b00010010;
		color_arr[165] = 8'b00010010;
		color_arr[166] = 8'b00010010;
		color_arr[167] = 8'b00010010;
		color_arr[168] = 8'b00010010;
		color_arr[169] = 8'b00010010;
		color_arr[170] = 8'b00010010;
		color_arr[171] = 8'b00010010;
		color_arr[172] = 8'b00010010;
		color_arr[173] = 8'b00010010;
		color_arr[174] = 8'b00010010;
		color_arr[175] = 8'b00010010;
		color_arr[176] = 8'b00010010;
		color_arr[177] = 8'b00010010;
		color_arr[178] = 8'b00010010;
		color_arr[179] = 8'b00010010;
		color_arr[180] = 8'b00010010;
		color_arr[181] = 8'b00010010;
		color_arr[182] = 8'b00010010;
		color_arr[183] = 8'b00010010;
		color_arr[184] = 8'b00010010;
		color_arr[185] = 8'b00010010;
		color_arr[186] = 8'b00010010;
		color_arr[187] = 8'b00000000;
		color_arr[188] = 8'b00000000;
		color_arr[189] = 8'b00000000;
		color_arr[190] = 8'b00000000;
		color_arr[191] = 8'b00000000;
		color_arr[192] = 8'b00000000;
		color_arr[193] = 8'b00000000;
		color_arr[194] = 8'b00000000;
		color_arr[195] = 8'b00000000;
		color_arr[196] = 8'b00000000;
		color_arr[197] = 8'b00000000;
		color_arr[198] = 8'b00000000;
		color_arr[199] = 8'b00000000;
		color_arr[200] = 8'b00000000;
		color_arr[201] = 8'b00010010;
		color_arr[202] = 8'b00010010;
		color_arr[203] = 8'b00010010;
		color_arr[204] = 8'b00010010;
		color_arr[205] = 8'b00000000;
		color_arr[206] = 8'b00000000;
		color_arr[207] = 8'b00000000;
		color_arr[208] = 8'b00000000;
		color_arr[209] = 8'b00000000;
		color_arr[210] = 8'b00000000;
		color_arr[211] = 8'b00000000;
		color_arr[212] = 8'b00010010;
		color_arr[213] = 8'b00010010;
		color_arr[214] = 8'b00010010;
		color_arr[215] = 8'b00010010;
		color_arr[216] = 8'b00010010;
		color_arr[217] = 8'b00010010;
		color_arr[218] = 8'b00010010;
		color_arr[219] = 8'b00010010;
		color_arr[220] = 8'b00010010;
		color_arr[221] = 8'b00010010;
		color_arr[222] = 8'b00010010;
		color_arr[223] = 8'b00010010;
		color_arr[224] = 8'b00010010;
		color_arr[225] = 8'b00010010;
		color_arr[226] = 8'b00010010;
		color_arr[227] = 8'b00010010;
		color_arr[228] = 8'b00010010;
		color_arr[229] = 8'b00010010;
		color_arr[230] = 8'b00010010;
		color_arr[231] = 8'b00010010;
		color_arr[232] = 8'b00010010;
		color_arr[233] = 8'b00010010;
		color_arr[234] = 8'b00010010;
		color_arr[235] = 8'b00010010;
		color_arr[236] = 8'b00010010;
		color_arr[237] = 8'b00010010;
		color_arr[238] = 8'b00010010;
		color_arr[239] = 8'b00010010;
		color_arr[240] = 8'b00010010;
		color_arr[241] = 8'b00010010;
		color_arr[242] = 8'b00010010;
		color_arr[243] = 8'b00010010;
		color_arr[244] = 8'b00010010;
		color_arr[245] = 8'b00010010;
		color_arr[246] = 8'b00010010;
		color_arr[247] = 8'b00010010;
		color_arr[248] = 8'b00010010;
		color_arr[249] = 8'b00010010;
		color_arr[250] = 8'b00010010;
		color_arr[251] = 8'b00010010;
		color_arr[252] = 8'b00010010;
		color_arr[253] = 8'b00010010;
		color_arr[254] = 8'b00010010;
		color_arr[255] = 8'b00010010;
		color_arr[256] = 8'b00010010;
		color_arr[257] = 8'b00010010;
		color_arr[258] = 8'b00010010;
		color_arr[259] = 8'b00010010;
		color_arr[260] = 8'b00010010;
		color_arr[261] = 8'b00010010;
		color_arr[262] = 8'b00010010;
		color_arr[263] = 8'b00010010;
		color_arr[264] = 8'b00010010;
		color_arr[265] = 8'b00010010;
		color_arr[266] = 8'b00010010;
		color_arr[267] = 8'b00010010;
		color_arr[268] = 8'b00010010;
		color_arr[269] = 8'b00010010;
		color_arr[270] = 8'b00010010;
		color_arr[271] = 8'b00010010;
		color_arr[272] = 8'b00010010;
		color_arr[273] = 8'b00010010;
		color_arr[274] = 8'b00010010;
		color_arr[275] = 8'b00010010;
		color_arr[276] = 8'b00010010;
		color_arr[277] = 8'b00010010;
		color_arr[278] = 8'b00010010;
		color_arr[279] = 8'b00010010;
		color_arr[280] = 8'b00010010;
		color_arr[281] = 8'b00010010;
		color_arr[282] = 8'b00010010;
		color_arr[283] = 8'b00010010;
		color_arr[284] = 8'b00010010;
		color_arr[285] = 8'b00010010;
		color_arr[286] = 8'b00010010;
		color_arr[287] = 8'b00010010;
		color_arr[288] = 8'b00010010;
		color_arr[289] = 8'b00010010;
		color_arr[290] = 8'b00010010;
		color_arr[291] = 8'b00010010;
		color_arr[292] = 8'b00010010;
		color_arr[293] = 8'b00010010;
		color_arr[294] = 8'b00010010;
		color_arr[295] = 8'b00010010;
		color_arr[296] = 8'b00010010;
		color_arr[297] = 8'b00010010;
		color_arr[298] = 8'b00010010;
		color_arr[299] = 8'b00010010;
		color_arr[300] = 8'b00010010;
		color_arr[301] = 8'b00010010;
		color_arr[302] = 8'b00010010;
		color_arr[303] = 8'b00010010;
		color_arr[304] = 8'b00010010;
		color_arr[305] = 8'b00010010;
		color_arr[306] = 8'b00010010;
		color_arr[307] = 8'b00010010;
		color_arr[308] = 8'b00010010;
		color_arr[309] = 8'b00010010;
		color_arr[310] = 8'b00010010;
		color_arr[311] = 8'b00010010;
		color_arr[312] = 8'b00000000;
		color_arr[313] = 8'b00000000;
		color_arr[314] = 8'b00000000;
		color_arr[315] = 8'b00000000;
		color_arr[316] = 8'b00000000;
		color_arr[317] = 8'b00000000;
		color_arr[318] = 8'b00000000;
		color_arr[319] = 8'b00000000;
		color_arr[320] = 8'b00000000;
		color_arr[321] = 8'b00010010;
		color_arr[322] = 8'b00010010;
		color_arr[323] = 8'b00010010;
		color_arr[324] = 8'b00010010;
		color_arr[325] = 8'b00010010;
		color_arr[326] = 8'b00010010;
		color_arr[327] = 8'b00010010;
		color_arr[328] = 8'b00010010;
		color_arr[329] = 8'b00010010;
		color_arr[330] = 8'b00010010;
		color_arr[331] = 8'b00010010;
		color_arr[332] = 8'b00010010;
		color_arr[333] = 8'b00010010;
		color_arr[334] = 8'b00010010;
		color_arr[335] = 8'b00010010;
		color_arr[336] = 8'b00000000;
		color_arr[337] = 8'b00000000;
		color_arr[338] = 8'b00000000;
		color_arr[339] = 8'b00000000;
		color_arr[340] = 8'b00000000;
		color_arr[341] = 8'b00000000;
		color_arr[342] = 8'b00010010;
		color_arr[343] = 8'b00010010;
		color_arr[344] = 8'b00010010;
		color_arr[345] = 8'b00010010;
		color_arr[346] = 8'b00010010;
		color_arr[347] = 8'b00010010;
		color_arr[348] = 8'b00010010;
		color_arr[349] = 8'b00010010;
		color_arr[350] = 8'b00010010;
		color_arr[351] = 8'b00010010;
		color_arr[352] = 8'b00010010;
		color_arr[353] = 8'b00010010;
		color_arr[354] = 8'b00010010;
		color_arr[355] = 8'b00010010;
		color_arr[356] = 8'b00010010;
		color_arr[357] = 8'b00010010;
		color_arr[358] = 8'b00010010;
		color_arr[359] = 8'b00010010;
		color_arr[360] = 8'b00010010;
		color_arr[361] = 8'b00010010;
		color_arr[362] = 8'b00010010;
		color_arr[363] = 8'b00010010;
		color_arr[364] = 8'b00010010;
		color_arr[365] = 8'b00010010;
		color_arr[366] = 8'b00010010;
		color_arr[367] = 8'b00010010;
		color_arr[368] = 8'b00010010;
		color_arr[369] = 8'b00010010;
		color_arr[370] = 8'b00010010;
		color_arr[371] = 8'b00010010;
		color_arr[372] = 8'b00010010;
		color_arr[373] = 8'b00010010;
		color_arr[374] = 8'b00010010;
		color_arr[375] = 8'b00010010;
		color_arr[376] = 8'b00010010;
		color_arr[377] = 8'b00010010;
		color_arr[378] = 8'b00010010;
		color_arr[379] = 8'b00010010;
		color_arr[380] = 8'b00010010;
		color_arr[381] = 8'b00010010;
		color_arr[382] = 8'b00010010;
		color_arr[383] = 8'b00010010;
		color_arr[384] = 8'b00010010;
		color_arr[385] = 8'b00010010;
		color_arr[386] = 8'b00010010;
		color_arr[387] = 8'b00010010;
		color_arr[388] = 8'b00010010;
		color_arr[389] = 8'b00010010;
		color_arr[390] = 8'b00010010;
		color_arr[391] = 8'b00010010;
		color_arr[392] = 8'b00010010;
		color_arr[393] = 8'b00010010;
		color_arr[394] = 8'b00010010;
		color_arr[395] = 8'b00010010;
		color_arr[396] = 8'b00010010;
		color_arr[397] = 8'b00010010;
		color_arr[398] = 8'b00010010;
		color_arr[399] = 8'b00010010;
		color_arr[400] = 8'b00010010;
		color_arr[401] = 8'b00010010;
		color_arr[402] = 8'b00010010;
		color_arr[403] = 8'b00010010;
		color_arr[404] = 8'b00010010;
		color_arr[405] = 8'b00010010;
		color_arr[406] = 8'b00010010;
		color_arr[407] = 8'b00010010;
		color_arr[408] = 8'b00010010;
		color_arr[409] = 8'b00010010;
		color_arr[410] = 8'b00010010;
		color_arr[411] = 8'b00010010;
		color_arr[412] = 8'b00010010;
		color_arr[413] = 8'b00010010;
		color_arr[414] = 8'b00010010;
		color_arr[415] = 8'b00010010;
		color_arr[416] = 8'b00010010;
		color_arr[417] = 8'b00010010;
		color_arr[418] = 8'b00010010;
		color_arr[419] = 8'b00010010;
		color_arr[420] = 8'b00010010;
		color_arr[421] = 8'b00010010;
		color_arr[422] = 8'b00010010;
		color_arr[423] = 8'b00010010;
		color_arr[424] = 8'b00010010;
		color_arr[425] = 8'b00010010;
		color_arr[426] = 8'b00010010;
		color_arr[427] = 8'b00010010;
		color_arr[428] = 8'b00010010;
		color_arr[429] = 8'b00010010;
		color_arr[430] = 8'b00010010;
		color_arr[431] = 8'b00010010;
		color_arr[432] = 8'b00010010;
		color_arr[433] = 8'b00010010;
		color_arr[434] = 8'b00010010;
		color_arr[435] = 8'b00010010;
		color_arr[436] = 8'b00010010;
		color_arr[437] = 8'b00010010;
		color_arr[438] = 8'b00000000;
		color_arr[439] = 8'b00000000;
		color_arr[440] = 8'b00000000;
		color_arr[441] = 8'b00000000;
		color_arr[442] = 8'b00000000;
		color_arr[443] = 8'b00000000;
		color_arr[444] = 8'b00010010;
		color_arr[445] = 8'b00010010;
		color_arr[446] = 8'b00010010;
		color_arr[447] = 8'b00010010;
		color_arr[448] = 8'b00010010;
		color_arr[449] = 8'b00010010;
		color_arr[450] = 8'b00010010;
		color_arr[451] = 8'b00010010;
		color_arr[452] = 8'b00010010;
		color_arr[453] = 8'b00010010;
		color_arr[454] = 8'b00010010;
		color_arr[455] = 8'b00010010;
		color_arr[456] = 8'b00010010;
		color_arr[457] = 8'b00010010;
		color_arr[458] = 8'b00010010;
		color_arr[459] = 8'b00010010;
		color_arr[460] = 8'b00010010;
		color_arr[461] = 8'b00010010;
		color_arr[462] = 8'b00010010;
		color_arr[463] = 8'b00010010;
		color_arr[464] = 8'b00010010;
		color_arr[465] = 8'b00010010;
		color_arr[466] = 8'b00010010;
		color_arr[467] = 8'b00000000;
		color_arr[468] = 8'b00000000;
		color_arr[469] = 8'b00000000;
		color_arr[470] = 8'b00000000;
		color_arr[471] = 8'b00000000;
		color_arr[472] = 8'b00010010;
		color_arr[473] = 8'b00010010;
		color_arr[474] = 8'b00010010;
		color_arr[475] = 8'b00010010;
		color_arr[476] = 8'b00010010;
		color_arr[477] = 8'b00010010;
		color_arr[478] = 8'b00010010;
		color_arr[479] = 8'b00010010;
		color_arr[480] = 8'b00010010;
		color_arr[481] = 8'b00010010;
		color_arr[482] = 8'b00010010;
		color_arr[483] = 8'b00010010;
		color_arr[484] = 8'b00010010;
		color_arr[485] = 8'b00010010;
		color_arr[486] = 8'b00010010;
		color_arr[487] = 8'b00010010;
		color_arr[488] = 8'b00010010;
		color_arr[489] = 8'b00010010;
		color_arr[490] = 8'b00010010;
		color_arr[491] = 8'b00010010;
		color_arr[492] = 8'b00010010;
		color_arr[493] = 8'b00010010;
		color_arr[494] = 8'b00010010;
		color_arr[495] = 8'b00010010;
		color_arr[496] = 8'b00010010;
		color_arr[497] = 8'b00010010;
		color_arr[498] = 8'b00010010;
		color_arr[499] = 8'b00010010;
		color_arr[500] = 8'b00010010;
		color_arr[501] = 8'b00010010;
		color_arr[502] = 8'b00010010;
		color_arr[503] = 8'b00010010;
		color_arr[504] = 8'b00010010;
		color_arr[505] = 8'b00010010;
		color_arr[506] = 8'b00010010;
		color_arr[507] = 8'b00010010;
		color_arr[508] = 8'b00010010;
		color_arr[509] = 8'b00010010;
		color_arr[510] = 8'b00010010;
		color_arr[511] = 8'b00010010;
		color_arr[512] = 8'b00010010;
		color_arr[513] = 8'b00010010;
		color_arr[514] = 8'b00010010;
		color_arr[515] = 8'b00010010;
		color_arr[516] = 8'b00010010;
		color_arr[517] = 8'b00010010;
		color_arr[518] = 8'b00010010;
		color_arr[519] = 8'b00010010;
		color_arr[520] = 8'b00010010;
		color_arr[521] = 8'b00010010;
		color_arr[522] = 8'b00010010;
		color_arr[523] = 8'b00010010;
		color_arr[524] = 8'b00010010;
		color_arr[525] = 8'b00010010;
		color_arr[526] = 8'b00010010;
		color_arr[527] = 8'b00010010;
		color_arr[528] = 8'b00010010;
		color_arr[529] = 8'b00010010;
		color_arr[530] = 8'b00010010;
		color_arr[531] = 8'b00010010;
		color_arr[532] = 8'b00010010;
		color_arr[533] = 8'b00010010;
		color_arr[534] = 8'b00010010;
		color_arr[535] = 8'b00010010;
		color_arr[536] = 8'b00010010;
		color_arr[537] = 8'b00010010;
		color_arr[538] = 8'b00010010;
		color_arr[539] = 8'b00010010;
		color_arr[540] = 8'b00010010;
		color_arr[541] = 8'b00010010;
		color_arr[542] = 8'b00010010;
		color_arr[543] = 8'b00010010;
		color_arr[544] = 8'b00010010;
		color_arr[545] = 8'b00010010;
		color_arr[546] = 8'b00010010;
		color_arr[547] = 8'b00010010;
		color_arr[548] = 8'b00010010;
		color_arr[549] = 8'b00010010;
		color_arr[550] = 8'b00010010;
		color_arr[551] = 8'b00010010;
		color_arr[552] = 8'b00010010;
		color_arr[553] = 8'b00010010;
		color_arr[554] = 8'b00010010;
		color_arr[555] = 8'b00010010;
		color_arr[556] = 8'b00010010;
		color_arr[557] = 8'b00010010;
		color_arr[558] = 8'b00010010;
		color_arr[559] = 8'b00010010;
		color_arr[560] = 8'b00010010;
		color_arr[561] = 8'b00010010;
		color_arr[562] = 8'b00010010;
		color_arr[563] = 8'b00010010;
		color_arr[564] = 8'b00000000;
		color_arr[565] = 8'b00000000;
		color_arr[566] = 8'b00000000;
		color_arr[567] = 8'b00000000;
		color_arr[568] = 8'b00000000;
		color_arr[569] = 8'b00010010;
		color_arr[570] = 8'b00010010;
		color_arr[571] = 8'b00010010;
		color_arr[572] = 8'b00010010;
		color_arr[573] = 8'b00010010;
		color_arr[574] = 8'b00010010;
		color_arr[575] = 8'b00010010;
		color_arr[576] = 8'b00010010;
		color_arr[577] = 8'b00010010;
		color_arr[578] = 8'b00010010;
		color_arr[579] = 8'b00010010;
		color_arr[580] = 8'b00010010;
		color_arr[581] = 8'b00010010;
		color_arr[582] = 8'b00010010;
		color_arr[583] = 8'b00010010;
		color_arr[584] = 8'b00010010;
		color_arr[585] = 8'b00010010;
		color_arr[586] = 8'b00010010;
		color_arr[587] = 8'b00010010;
		color_arr[588] = 8'b00010010;
		color_arr[589] = 8'b00010010;
		color_arr[590] = 8'b00010010;
		color_arr[591] = 8'b00010010;
		color_arr[592] = 8'b00010010;
		color_arr[593] = 8'b00010010;
		color_arr[594] = 8'b00010010;
		color_arr[595] = 8'b00010010;
		color_arr[596] = 8'b00010010;
		color_arr[597] = 8'b00000000;
		color_arr[598] = 8'b00000000;
		color_arr[599] = 8'b00000000;
		color_arr[600] = 8'b00000000;
		color_arr[601] = 8'b00010010;
		color_arr[602] = 8'b00010010;
		color_arr[603] = 8'b00010010;
		color_arr[604] = 8'b00010010;
		color_arr[605] = 8'b00010010;
		color_arr[606] = 8'b00010010;
		color_arr[607] = 8'b00010010;
		color_arr[608] = 8'b00010010;
		color_arr[609] = 8'b00010010;
		color_arr[610] = 8'b00010010;
		color_arr[611] = 8'b00010010;
		color_arr[612] = 8'b00010010;
		color_arr[613] = 8'b00010010;
		color_arr[614] = 8'b00010010;
		color_arr[615] = 8'b00010010;
		color_arr[616] = 8'b00010010;
		color_arr[617] = 8'b00010010;
		color_arr[618] = 8'b00010010;
		color_arr[619] = 8'b00010010;
		color_arr[620] = 8'b00010010;
		color_arr[621] = 8'b00010010;
		color_arr[622] = 8'b00010010;
		color_arr[623] = 8'b00010010;
		color_arr[624] = 8'b00010010;
		color_arr[625] = 8'b00010010;
		color_arr[626] = 8'b00010010;
		color_arr[627] = 8'b00010010;
		color_arr[628] = 8'b00010010;
		color_arr[629] = 8'b00010010;
		color_arr[630] = 8'b00010010;
		color_arr[631] = 8'b00010010;
		color_arr[632] = 8'b00010010;
		color_arr[633] = 8'b00010010;
		color_arr[634] = 8'b00010010;
		color_arr[635] = 8'b00010010;
		color_arr[636] = 8'b00010010;
		color_arr[637] = 8'b00010010;
		color_arr[638] = 8'b00010010;
		color_arr[639] = 8'b00010010;
		color_arr[640] = 8'b00010010;
		color_arr[641] = 8'b00010010;
		color_arr[642] = 8'b00010010;
		color_arr[643] = 8'b00010010;
		color_arr[644] = 8'b00010010;
		color_arr[645] = 8'b00010010;
		color_arr[646] = 8'b00010010;
		color_arr[647] = 8'b00010010;
		color_arr[648] = 8'b00010010;
		color_arr[649] = 8'b00010010;
		color_arr[650] = 8'b00010010;
		color_arr[651] = 8'b00010010;
		color_arr[652] = 8'b00010010;
		color_arr[653] = 8'b00010010;
		color_arr[654] = 8'b00010010;
		color_arr[655] = 8'b00010010;
		color_arr[656] = 8'b00010010;
		color_arr[657] = 8'b00010010;
		color_arr[658] = 8'b00010010;
		color_arr[659] = 8'b00010010;
		color_arr[660] = 8'b00010010;
		color_arr[661] = 8'b00010010;
		color_arr[662] = 8'b00010010;
		color_arr[663] = 8'b00010010;
		color_arr[664] = 8'b00010010;
		color_arr[665] = 8'b00010010;
		color_arr[666] = 8'b00010010;
		color_arr[667] = 8'b00010010;
		color_arr[668] = 8'b00010010;
		color_arr[669] = 8'b00010010;
		color_arr[670] = 8'b00010010;
		color_arr[671] = 8'b00010010;
		color_arr[672] = 8'b00010010;
		color_arr[673] = 8'b00010010;
		color_arr[674] = 8'b00010010;
		color_arr[675] = 8'b00010010;
		color_arr[676] = 8'b00010010;
		color_arr[677] = 8'b00010010;
		color_arr[678] = 8'b00010010;
		color_arr[679] = 8'b00010010;
		color_arr[680] = 8'b00010010;
		color_arr[681] = 8'b00010010;
		color_arr[682] = 8'b00010010;
		color_arr[683] = 8'b00010010;
		color_arr[684] = 8'b00010010;
		color_arr[685] = 8'b00010010;
		color_arr[686] = 8'b00010010;
		color_arr[687] = 8'b00010010;
		color_arr[688] = 8'b00010010;
		color_arr[689] = 8'b00010010;
		color_arr[690] = 8'b00000000;
		color_arr[691] = 8'b00000000;
		color_arr[692] = 8'b00000000;
		color_arr[693] = 8'b00000000;
		color_arr[694] = 8'b00000000;
		color_arr[695] = 8'b00010010;
		color_arr[696] = 8'b00010010;
		color_arr[697] = 8'b00010010;
		color_arr[698] = 8'b00010010;
		color_arr[699] = 8'b00010010;
		color_arr[700] = 8'b00010010;
		color_arr[701] = 8'b00010010;
		color_arr[702] = 8'b00010010;
		color_arr[703] = 8'b00010010;
		color_arr[704] = 8'b00010010;
		color_arr[705] = 8'b00010010;
		color_arr[706] = 8'b00010010;
		color_arr[707] = 8'b00010010;
		color_arr[708] = 8'b00010010;
		color_arr[709] = 8'b00010010;
		color_arr[710] = 8'b00010010;
		color_arr[711] = 8'b00010010;
		color_arr[712] = 8'b00010010;
		color_arr[713] = 8'b00010010;
		color_arr[714] = 8'b00010010;
		color_arr[715] = 8'b00010010;
		color_arr[716] = 8'b00010010;
		color_arr[717] = 8'b00010010;
		color_arr[718] = 8'b00010010;
		color_arr[719] = 8'b00010010;
		color_arr[720] = 8'b00010010;
		color_arr[721] = 8'b00010010;
		color_arr[722] = 8'b00010010;
		color_arr[723] = 8'b00010010;
		color_arr[724] = 8'b00010010;
		color_arr[725] = 8'b00010010;
		color_arr[726] = 8'b00010010;
		color_arr[727] = 8'b00000000;
		color_arr[728] = 8'b00000000;
		color_arr[729] = 8'b00000000;
		color_arr[730] = 8'b00000000;
		color_arr[731] = 8'b00010010;
		color_arr[732] = 8'b00010010;
		color_arr[733] = 8'b00010010;
		color_arr[734] = 8'b00010010;
		color_arr[735] = 8'b00010010;
		color_arr[736] = 8'b00010010;
		color_arr[737] = 8'b00010010;
		color_arr[738] = 8'b00010010;
		color_arr[739] = 8'b00010010;
		color_arr[740] = 8'b00010010;
		color_arr[741] = 8'b00010010;
		color_arr[742] = 8'b00010010;
		color_arr[743] = 8'b00010010;
		color_arr[744] = 8'b00010010;
		color_arr[745] = 8'b00010010;
		color_arr[746] = 8'b00010010;
		color_arr[747] = 8'b00010010;
		color_arr[748] = 8'b00010010;
		color_arr[749] = 8'b00010010;
		color_arr[750] = 8'b00010010;
		color_arr[751] = 8'b00010010;
		color_arr[752] = 8'b00010010;
		color_arr[753] = 8'b00010010;
		color_arr[754] = 8'b00010010;
		color_arr[755] = 8'b00010010;
		color_arr[756] = 8'b00010010;
		color_arr[757] = 8'b00010010;
		color_arr[758] = 8'b00010010;
		color_arr[759] = 8'b00010010;
		color_arr[760] = 8'b00010010;
		color_arr[761] = 8'b00010010;
		color_arr[762] = 8'b00010010;
		color_arr[763] = 8'b00010010;
		color_arr[764] = 8'b00010010;
		color_arr[765] = 8'b00010010;
		color_arr[766] = 8'b00010010;
		color_arr[767] = 8'b00010010;
		color_arr[768] = 8'b00010010;
		color_arr[769] = 8'b00010010;
		color_arr[770] = 8'b00010010;
		color_arr[771] = 8'b00010010;
		color_arr[772] = 8'b00010010;
		color_arr[773] = 8'b00010010;
		color_arr[774] = 8'b00010010;
		color_arr[775] = 8'b00010010;
		color_arr[776] = 8'b00010010;
		color_arr[777] = 8'b00010010;
		color_arr[778] = 8'b00010010;
		color_arr[779] = 8'b00010010;
		color_arr[780] = 8'b00010010;
		color_arr[781] = 8'b00010010;
		color_arr[782] = 8'b00010010;
		color_arr[783] = 8'b00010010;
		color_arr[784] = 8'b00010010;
		color_arr[785] = 8'b00010010;
		color_arr[786] = 8'b00010010;
		color_arr[787] = 8'b00010010;
		color_arr[788] = 8'b00010010;
		color_arr[789] = 8'b00010010;
		color_arr[790] = 8'b00010010;
		color_arr[791] = 8'b00010010;
		color_arr[792] = 8'b00010010;
		color_arr[793] = 8'b00010010;
		color_arr[794] = 8'b00010010;
		color_arr[795] = 8'b00010010;
		color_arr[796] = 8'b00010010;
		color_arr[797] = 8'b00010010;
		color_arr[798] = 8'b00010010;
		color_arr[799] = 8'b00010010;
		color_arr[800] = 8'b00010010;
		color_arr[801] = 8'b00010010;
		color_arr[802] = 8'b00010010;
		color_arr[803] = 8'b00010010;
		color_arr[804] = 8'b00010010;
		color_arr[805] = 8'b00010010;
		color_arr[806] = 8'b00010010;
		color_arr[807] = 8'b00010010;
		color_arr[808] = 8'b00010010;
		color_arr[809] = 8'b00010010;
		color_arr[810] = 8'b00010010;
		color_arr[811] = 8'b00010010;
		color_arr[812] = 8'b00010010;
		color_arr[813] = 8'b00010010;
		color_arr[814] = 8'b00010010;
		color_arr[815] = 8'b00010010;
		color_arr[816] = 8'b00000000;
		color_arr[817] = 8'b00000000;
		color_arr[818] = 8'b00000000;
		color_arr[819] = 8'b00000000;
		color_arr[820] = 8'b00000000;
		color_arr[821] = 8'b00010010;
		color_arr[822] = 8'b00010010;
		color_arr[823] = 8'b00010010;
		color_arr[824] = 8'b00010010;
		color_arr[825] = 8'b00010010;
		color_arr[826] = 8'b00010010;
		color_arr[827] = 8'b00010010;
		color_arr[828] = 8'b00010010;
		color_arr[829] = 8'b00010010;
		color_arr[830] = 8'b00010010;
		color_arr[831] = 8'b00010010;
		color_arr[832] = 8'b00010010;
		color_arr[833] = 8'b00010010;
		color_arr[834] = 8'b00010010;
		color_arr[835] = 8'b00010010;
		color_arr[836] = 8'b00010010;
		color_arr[837] = 8'b00010010;
		color_arr[838] = 8'b00010010;
		color_arr[839] = 8'b00010010;
		color_arr[840] = 8'b00010010;
		color_arr[841] = 8'b00010010;
		color_arr[842] = 8'b00010010;
		color_arr[843] = 8'b00010010;
		color_arr[844] = 8'b00010010;
		color_arr[845] = 8'b00010010;
		color_arr[846] = 8'b00010010;
		color_arr[847] = 8'b00010010;
		color_arr[848] = 8'b00100000;
		color_arr[849] = 8'b00100000;
		color_arr[850] = 8'b00100000;
		color_arr[851] = 8'b00100000;
		color_arr[852] = 8'b00100000;
		color_arr[853] = 8'b00100000;
		color_arr[854] = 8'b00100000;
		color_arr[855] = 8'b00100000;
		color_arr[856] = 8'b00000000;
		color_arr[857] = 8'b00000000;
		color_arr[858] = 8'b00000000;
		color_arr[859] = 8'b00000000;
		color_arr[860] = 8'b00000000;
		color_arr[861] = 8'b00000000;
		color_arr[862] = 8'b00000000;
		color_arr[863] = 8'b00000000;
		color_arr[864] = 8'b00000000;
		color_arr[865] = 8'b00000000;
		color_arr[866] = 8'b00000000;
		color_arr[867] = 8'b00000000;
		color_arr[868] = 8'b00000000;
		color_arr[869] = 8'b00100000;
		color_arr[870] = 8'b00100000;
		color_arr[871] = 8'b00100000;
		color_arr[872] = 8'b00100000;
		color_arr[873] = 8'b00100000;
		color_arr[874] = 8'b00100000;
		color_arr[875] = 8'b00100000;
		color_arr[876] = 8'b00100000;
		color_arr[877] = 8'b00100000;
		color_arr[878] = 8'b00100000;
		color_arr[879] = 8'b00100000;
		color_arr[880] = 8'b00100000;
		color_arr[881] = 8'b00100000;
		color_arr[882] = 8'b00100000;
		color_arr[883] = 8'b00100000;
		color_arr[884] = 8'b00100000;
		color_arr[885] = 8'b00100000;
		color_arr[886] = 8'b00100000;
		color_arr[887] = 8'b00100000;
		color_arr[888] = 8'b00100000;
		color_arr[889] = 8'b00100000;
		color_arr[890] = 8'b00100000;
		color_arr[891] = 8'b00100000;
		color_arr[892] = 8'b00100000;
		color_arr[893] = 8'b00010010;
		color_arr[894] = 8'b00010010;
		color_arr[895] = 8'b00010010;
		color_arr[896] = 8'b00010010;
		color_arr[897] = 8'b00010010;
		color_arr[898] = 8'b00010010;
		color_arr[899] = 8'b00010010;
		color_arr[900] = 8'b00010010;
		color_arr[901] = 8'b00010010;
		color_arr[902] = 8'b00010010;
		color_arr[903] = 8'b00010010;
		color_arr[904] = 8'b00010010;
		color_arr[905] = 8'b00010010;
		color_arr[906] = 8'b00010010;
		color_arr[907] = 8'b00010010;
		color_arr[908] = 8'b00010010;
		color_arr[909] = 8'b00010010;
		color_arr[910] = 8'b00010010;
		color_arr[911] = 8'b00010010;
		color_arr[912] = 8'b00010010;
		color_arr[913] = 8'b00010010;
		color_arr[914] = 8'b00010010;
		color_arr[915] = 8'b00010010;
		color_arr[916] = 8'b00010010;
		color_arr[917] = 8'b00010010;
		color_arr[918] = 8'b00010010;
		color_arr[919] = 8'b00010010;
		color_arr[920] = 8'b00010010;
		color_arr[921] = 8'b00010010;
		color_arr[922] = 8'b00010010;
		color_arr[923] = 8'b00010010;
		color_arr[924] = 8'b00010010;
		color_arr[925] = 8'b00010010;
		color_arr[926] = 8'b00010010;
		color_arr[927] = 8'b00010010;
		color_arr[928] = 8'b00010010;
		color_arr[929] = 8'b00010010;
		color_arr[930] = 8'b00010010;
		color_arr[931] = 8'b00010010;
		color_arr[932] = 8'b00010010;
		color_arr[933] = 8'b00010010;
		color_arr[934] = 8'b00010010;
		color_arr[935] = 8'b00010010;
		color_arr[936] = 8'b00010010;
		color_arr[937] = 8'b00010010;
		color_arr[938] = 8'b00010010;
		color_arr[939] = 8'b00010010;
		color_arr[940] = 8'b00010010;
		color_arr[941] = 8'b00010010;
		color_arr[942] = 8'b00000000;
		color_arr[943] = 8'b00000000;
		color_arr[944] = 8'b00000000;
		color_arr[945] = 8'b00000000;
		color_arr[946] = 8'b00000000;
		color_arr[947] = 8'b00010010;
		color_arr[948] = 8'b00010010;
		color_arr[949] = 8'b00010010;
		color_arr[950] = 8'b00010010;
		color_arr[951] = 8'b00010010;
		color_arr[952] = 8'b00010010;
		color_arr[953] = 8'b00010010;
		color_arr[954] = 8'b00010010;
		color_arr[955] = 8'b00010010;
		color_arr[956] = 8'b00010010;
		color_arr[957] = 8'b00010010;
		color_arr[958] = 8'b00010010;
		color_arr[959] = 8'b00010010;
		color_arr[960] = 8'b00010010;
		color_arr[961] = 8'b00010010;
		color_arr[962] = 8'b00010010;
		color_arr[963] = 8'b00010010;
		color_arr[964] = 8'b00010010;
		color_arr[965] = 8'b00010010;
		color_arr[966] = 8'b00010010;
		color_arr[967] = 8'b00010010;
		color_arr[968] = 8'b00010010;
		color_arr[969] = 8'b00010010;
		color_arr[970] = 8'b00010010;
		color_arr[971] = 8'b00010010;
		color_arr[972] = 8'b00010010;
		color_arr[973] = 8'b00010010;
		color_arr[974] = 8'b00010010;
		color_arr[975] = 8'b00010010;
		color_arr[976] = 8'b00100000;
		color_arr[977] = 8'b00100000;
		color_arr[978] = 8'b00100000;
		color_arr[979] = 8'b00100000;
		color_arr[980] = 8'b00100000;
		color_arr[981] = 8'b00100000;
		color_arr[982] = 8'b00100000;
		color_arr[983] = 8'b00100000;
		color_arr[984] = 8'b00100000;
		color_arr[985] = 8'b00100000;
		color_arr[986] = 8'b00000000;
		color_arr[987] = 8'b00000000;
		color_arr[988] = 8'b00000000;
		color_arr[989] = 8'b00000000;
		color_arr[990] = 8'b00000000;
		color_arr[991] = 8'b00000000;
		color_arr[992] = 8'b00000000;
		color_arr[993] = 8'b00000000;
		color_arr[994] = 8'b00000000;
		color_arr[995] = 8'b00000000;
		color_arr[996] = 8'b00000000;
		color_arr[997] = 8'b00000000;
		color_arr[998] = 8'b00000000;
		color_arr[999] = 8'b00000000;
		color_arr[1000] = 8'b00000000;
		color_arr[1001] = 8'b00000000;
		color_arr[1002] = 8'b00100000;
		color_arr[1003] = 8'b00100000;
		color_arr[1004] = 8'b00100000;
		color_arr[1005] = 8'b00100000;
		color_arr[1006] = 8'b00100000;
		color_arr[1007] = 8'b00100000;
		color_arr[1008] = 8'b00100000;
		color_arr[1009] = 8'b00100000;
		color_arr[1010] = 8'b00100000;
		color_arr[1011] = 8'b00100000;
		color_arr[1012] = 8'b00100000;
		color_arr[1013] = 8'b00100000;
		color_arr[1014] = 8'b00100000;
		color_arr[1015] = 8'b00100000;
		color_arr[1016] = 8'b00100000;
		color_arr[1017] = 8'b00100000;
		color_arr[1018] = 8'b00100000;
		color_arr[1019] = 8'b00100000;
		color_arr[1020] = 8'b00100000;
		color_arr[1021] = 8'b00010010;
		color_arr[1022] = 8'b00010010;
		color_arr[1023] = 8'b00010010;
		color_arr[1024] = 8'b00010010;
		color_arr[1025] = 8'b00010010;
		color_arr[1026] = 8'b00010010;
		color_arr[1027] = 8'b00010010;
		color_arr[1028] = 8'b00010010;
		color_arr[1029] = 8'b00010010;
		color_arr[1030] = 8'b00010010;
		color_arr[1031] = 8'b00010010;
		color_arr[1032] = 8'b00000010;
		color_arr[1033] = 8'b00000010;
		color_arr[1034] = 8'b00000010;
		color_arr[1035] = 8'b00000010;
		color_arr[1036] = 8'b00000010;
		color_arr[1037] = 8'b00000010;
		color_arr[1038] = 8'b00000010;
		color_arr[1039] = 8'b00000010;
		color_arr[1040] = 8'b00000010;
		color_arr[1041] = 8'b00000010;
		color_arr[1042] = 8'b00000010;
		color_arr[1043] = 8'b00000010;
		color_arr[1044] = 8'b00000010;
		color_arr[1045] = 8'b00000010;
		color_arr[1046] = 8'b00000010;
		color_arr[1047] = 8'b00000010;
		color_arr[1048] = 8'b00000010;
		color_arr[1049] = 8'b00000010;
		color_arr[1050] = 8'b00000010;
		color_arr[1051] = 8'b00000010;
		color_arr[1052] = 8'b00000010;
		color_arr[1053] = 8'b00000010;
		color_arr[1054] = 8'b00000010;
		color_arr[1055] = 8'b00000010;
		color_arr[1056] = 8'b00000010;
		color_arr[1057] = 8'b00000010;
		color_arr[1058] = 8'b00000010;
		color_arr[1059] = 8'b00000010;
		color_arr[1060] = 8'b00000010;
		color_arr[1061] = 8'b00000010;
		color_arr[1062] = 8'b00010010;
		color_arr[1063] = 8'b00010010;
		color_arr[1064] = 8'b00010010;
		color_arr[1065] = 8'b00010010;
		color_arr[1066] = 8'b00010010;
		color_arr[1067] = 8'b00010010;
		color_arr[1068] = 8'b00000000;
		color_arr[1069] = 8'b00000000;
		color_arr[1070] = 8'b00000000;
		color_arr[1071] = 8'b00000000;
		color_arr[1072] = 8'b00000000;
		color_arr[1073] = 8'b00010010;
		color_arr[1074] = 8'b00010010;
		color_arr[1075] = 8'b00010010;
		color_arr[1076] = 8'b00010010;
		color_arr[1077] = 8'b00010010;
		color_arr[1078] = 8'b00010010;
		color_arr[1079] = 8'b00010010;
		color_arr[1080] = 8'b00010010;
		color_arr[1081] = 8'b00010010;
		color_arr[1082] = 8'b00010010;
		color_arr[1083] = 8'b00010010;
		color_arr[1084] = 8'b00010010;
		color_arr[1085] = 8'b00010010;
		color_arr[1086] = 8'b00010010;
		color_arr[1087] = 8'b00010010;
		color_arr[1088] = 8'b00010010;
		color_arr[1089] = 8'b00010010;
		color_arr[1090] = 8'b00010010;
		color_arr[1091] = 8'b00010010;
		color_arr[1092] = 8'b00010010;
		color_arr[1093] = 8'b00010010;
		color_arr[1094] = 8'b00010010;
		color_arr[1095] = 8'b00010010;
		color_arr[1096] = 8'b00010010;
		color_arr[1097] = 8'b00010010;
		color_arr[1098] = 8'b00010010;
		color_arr[1099] = 8'b00010010;
		color_arr[1100] = 8'b00010010;
		color_arr[1101] = 8'b00010010;
		color_arr[1102] = 8'b00010010;
		color_arr[1103] = 8'b00010010;
		color_arr[1104] = 8'b00100000;
		color_arr[1105] = 8'b00100000;
		color_arr[1106] = 8'b00100000;
		color_arr[1107] = 8'b00100000;
		color_arr[1108] = 8'b00100000;
		color_arr[1109] = 8'b00100000;
		color_arr[1110] = 8'b00100000;
		color_arr[1111] = 8'b00100000;
		color_arr[1112] = 8'b00100000;
		color_arr[1113] = 8'b00100000;
		color_arr[1114] = 8'b00100000;
		color_arr[1115] = 8'b00000000;
		color_arr[1116] = 8'b00000000;
		color_arr[1117] = 8'b00000000;
		color_arr[1118] = 8'b00100000;
		color_arr[1119] = 8'b00100000;
		color_arr[1120] = 8'b00100000;
		color_arr[1121] = 8'b00100000;
		color_arr[1122] = 8'b00100000;
		color_arr[1123] = 8'b00100000;
		color_arr[1124] = 8'b00000000;
		color_arr[1125] = 8'b00000000;
		color_arr[1126] = 8'b00000000;
		color_arr[1127] = 8'b00000000;
		color_arr[1128] = 8'b00000000;
		color_arr[1129] = 8'b00000000;
		color_arr[1130] = 8'b00000000;
		color_arr[1131] = 8'b00000000;
		color_arr[1132] = 8'b00000000;
		color_arr[1133] = 8'b00100000;
		color_arr[1134] = 8'b00100000;
		color_arr[1135] = 8'b00100000;
		color_arr[1136] = 8'b00100000;
		color_arr[1137] = 8'b00100000;
		color_arr[1138] = 8'b00100000;
		color_arr[1139] = 8'b00100000;
		color_arr[1140] = 8'b00100000;
		color_arr[1141] = 8'b00100000;
		color_arr[1142] = 8'b00100000;
		color_arr[1143] = 8'b00100000;
		color_arr[1144] = 8'b00100000;
		color_arr[1145] = 8'b00100000;
		color_arr[1146] = 8'b00100000;
		color_arr[1147] = 8'b00100000;
		color_arr[1148] = 8'b00100000;
		color_arr[1149] = 8'b00010010;
		color_arr[1150] = 8'b00010010;
		color_arr[1151] = 8'b00010010;
		color_arr[1152] = 8'b00010010;
		color_arr[1153] = 8'b00010010;
		color_arr[1154] = 8'b00010010;
		color_arr[1155] = 8'b00010010;
		color_arr[1156] = 8'b00010010;
		color_arr[1157] = 8'b00010010;
		color_arr[1158] = 8'b00010010;
		color_arr[1159] = 8'b00010010;
		color_arr[1160] = 8'b00000010;
		color_arr[1161] = 8'b00000010;
		color_arr[1162] = 8'b00000010;
		color_arr[1163] = 8'b00000010;
		color_arr[1164] = 8'b00000010;
		color_arr[1165] = 8'b00000010;
		color_arr[1166] = 8'b00000010;
		color_arr[1167] = 8'b00000010;
		color_arr[1168] = 8'b00000010;
		color_arr[1169] = 8'b00000010;
		color_arr[1170] = 8'b00000010;
		color_arr[1171] = 8'b00000010;
		color_arr[1172] = 8'b00000010;
		color_arr[1173] = 8'b00000010;
		color_arr[1174] = 8'b00000010;
		color_arr[1175] = 8'b00000010;
		color_arr[1176] = 8'b00000010;
		color_arr[1177] = 8'b00000010;
		color_arr[1178] = 8'b00000010;
		color_arr[1179] = 8'b00000010;
		color_arr[1180] = 8'b00000010;
		color_arr[1181] = 8'b00000010;
		color_arr[1182] = 8'b00000010;
		color_arr[1183] = 8'b00000010;
		color_arr[1184] = 8'b00000010;
		color_arr[1185] = 8'b00000010;
		color_arr[1186] = 8'b00000010;
		color_arr[1187] = 8'b00000010;
		color_arr[1188] = 8'b00000010;
		color_arr[1189] = 8'b00000010;
		color_arr[1190] = 8'b00010010;
		color_arr[1191] = 8'b00010010;
		color_arr[1192] = 8'b00010010;
		color_arr[1193] = 8'b00010010;
		color_arr[1194] = 8'b00010010;
		color_arr[1195] = 8'b00000000;
		color_arr[1196] = 8'b00000000;
		color_arr[1197] = 8'b00000000;
		color_arr[1198] = 8'b00000000;
		color_arr[1199] = 8'b00010010;
		color_arr[1200] = 8'b00010010;
		color_arr[1201] = 8'b00010010;
		color_arr[1202] = 8'b00010010;
		color_arr[1203] = 8'b00010010;
		color_arr[1204] = 8'b00010010;
		color_arr[1205] = 8'b00010010;
		color_arr[1206] = 8'b00010010;
		color_arr[1207] = 8'b00010010;
		color_arr[1208] = 8'b00010010;
		color_arr[1209] = 8'b00010010;
		color_arr[1210] = 8'b00010010;
		color_arr[1211] = 8'b00010010;
		color_arr[1212] = 8'b00010010;
		color_arr[1213] = 8'b00010010;
		color_arr[1214] = 8'b00010010;
		color_arr[1215] = 8'b00010010;
		color_arr[1216] = 8'b00010010;
		color_arr[1217] = 8'b00010010;
		color_arr[1218] = 8'b00010010;
		color_arr[1219] = 8'b00010010;
		color_arr[1220] = 8'b00010010;
		color_arr[1221] = 8'b00010010;
		color_arr[1222] = 8'b00010010;
		color_arr[1223] = 8'b00010010;
		color_arr[1224] = 8'b00010010;
		color_arr[1225] = 8'b00010010;
		color_arr[1226] = 8'b00010010;
		color_arr[1227] = 8'b00010010;
		color_arr[1228] = 8'b00010010;
		color_arr[1229] = 8'b00010010;
		color_arr[1230] = 8'b00010010;
		color_arr[1231] = 8'b00010010;
		color_arr[1232] = 8'b00100000;
		color_arr[1233] = 8'b00100000;
		color_arr[1234] = 8'b00100000;
		color_arr[1235] = 8'b00100000;
		color_arr[1236] = 8'b00100000;
		color_arr[1237] = 8'b00100000;
		color_arr[1238] = 8'b00100000;
		color_arr[1239] = 8'b00100000;
		color_arr[1240] = 8'b00100000;
		color_arr[1241] = 8'b00100000;
		color_arr[1242] = 8'b00100000;
		color_arr[1243] = 8'b00100000;
		color_arr[1244] = 8'b00000000;
		color_arr[1245] = 8'b00000000;
		color_arr[1246] = 8'b00100000;
		color_arr[1247] = 8'b00100000;
		color_arr[1248] = 8'b00100000;
		color_arr[1249] = 8'b00100000;
		color_arr[1250] = 8'b00100000;
		color_arr[1251] = 8'b00100000;
		color_arr[1252] = 8'b00100000;
		color_arr[1253] = 8'b00100000;
		color_arr[1254] = 8'b00100000;
		color_arr[1255] = 8'b00100000;
		color_arr[1256] = 8'b00100000;
		color_arr[1257] = 8'b00000000;
		color_arr[1258] = 8'b00000000;
		color_arr[1259] = 8'b00000000;
		color_arr[1260] = 8'b00000000;
		color_arr[1261] = 8'b00000000;
		color_arr[1262] = 8'b00100000;
		color_arr[1263] = 8'b00100000;
		color_arr[1264] = 8'b00100000;
		color_arr[1265] = 8'b00100000;
		color_arr[1266] = 8'b00100000;
		color_arr[1267] = 8'b00100000;
		color_arr[1268] = 8'b00100000;
		color_arr[1269] = 8'b00100000;
		color_arr[1270] = 8'b00100000;
		color_arr[1271] = 8'b00100000;
		color_arr[1272] = 8'b00100000;
		color_arr[1273] = 8'b00100000;
		color_arr[1274] = 8'b00100000;
		color_arr[1275] = 8'b00100000;
		color_arr[1276] = 8'b00100000;
		color_arr[1277] = 8'b00010010;
		color_arr[1278] = 8'b00010010;
		color_arr[1279] = 8'b00010010;
		color_arr[1280] = 8'b00010010;
		color_arr[1281] = 8'b00010010;
		color_arr[1282] = 8'b00010010;
		color_arr[1283] = 8'b00010010;
		color_arr[1284] = 8'b00010010;
		color_arr[1285] = 8'b00010010;
		color_arr[1286] = 8'b00010010;
		color_arr[1287] = 8'b00010010;
		color_arr[1288] = 8'b00000010;
		color_arr[1289] = 8'b00000010;
		color_arr[1290] = 8'b00000010;
		color_arr[1291] = 8'b00000010;
		color_arr[1292] = 8'b00000010;
		color_arr[1293] = 8'b00000010;
		color_arr[1294] = 8'b00000010;
		color_arr[1295] = 8'b00000010;
		color_arr[1296] = 8'b00000010;
		color_arr[1297] = 8'b00000010;
		color_arr[1298] = 8'b00000010;
		color_arr[1299] = 8'b00000010;
		color_arr[1300] = 8'b00000010;
		color_arr[1301] = 8'b00000010;
		color_arr[1302] = 8'b00000010;
		color_arr[1303] = 8'b00000010;
		color_arr[1304] = 8'b00000010;
		color_arr[1305] = 8'b00000010;
		color_arr[1306] = 8'b00000010;
		color_arr[1307] = 8'b00000010;
		color_arr[1308] = 8'b00000010;
		color_arr[1309] = 8'b00000010;
		color_arr[1310] = 8'b00000010;
		color_arr[1311] = 8'b00000010;
		color_arr[1312] = 8'b00000010;
		color_arr[1313] = 8'b00000010;
		color_arr[1314] = 8'b00000010;
		color_arr[1315] = 8'b00000010;
		color_arr[1316] = 8'b00000010;
		color_arr[1317] = 8'b00000010;
		color_arr[1318] = 8'b00010010;
		color_arr[1319] = 8'b00010010;
		color_arr[1320] = 8'b00010010;
		color_arr[1321] = 8'b00000000;
		color_arr[1322] = 8'b00000000;
		color_arr[1323] = 8'b00000000;
		color_arr[1324] = 8'b00000000;
		color_arr[1325] = 8'b00010010;
		color_arr[1326] = 8'b00010010;
		color_arr[1327] = 8'b00010010;
		color_arr[1328] = 8'b00010010;
		color_arr[1329] = 8'b00010010;
		color_arr[1330] = 8'b00010010;
		color_arr[1331] = 8'b00010010;
		color_arr[1332] = 8'b00010010;
		color_arr[1333] = 8'b00010010;
		color_arr[1334] = 8'b00010010;
		color_arr[1335] = 8'b00010010;
		color_arr[1336] = 8'b00010010;
		color_arr[1337] = 8'b00010010;
		color_arr[1338] = 8'b00010010;
		color_arr[1339] = 8'b00010010;
		color_arr[1340] = 8'b00010010;
		color_arr[1341] = 8'b00010010;
		color_arr[1342] = 8'b00010010;
		color_arr[1343] = 8'b00010010;
		color_arr[1344] = 8'b00010010;
		color_arr[1345] = 8'b00010010;
		color_arr[1346] = 8'b00010010;
		color_arr[1347] = 8'b00010010;
		color_arr[1348] = 8'b00010010;
		color_arr[1349] = 8'b00010010;
		color_arr[1350] = 8'b00010010;
		color_arr[1351] = 8'b00010010;
		color_arr[1352] = 8'b00010010;
		color_arr[1353] = 8'b00010010;
		color_arr[1354] = 8'b00010010;
		color_arr[1355] = 8'b00010010;
		color_arr[1356] = 8'b00010010;
		color_arr[1357] = 8'b00010010;
		color_arr[1358] = 8'b00010010;
		color_arr[1359] = 8'b00010010;
		color_arr[1360] = 8'b00100000;
		color_arr[1361] = 8'b00100000;
		color_arr[1362] = 8'b00100000;
		color_arr[1363] = 8'b00100000;
		color_arr[1364] = 8'b00100000;
		color_arr[1365] = 8'b00100000;
		color_arr[1366] = 8'b00100000;
		color_arr[1367] = 8'b00100000;
		color_arr[1368] = 8'b00100000;
		color_arr[1369] = 8'b00100000;
		color_arr[1370] = 8'b00100000;
		color_arr[1371] = 8'b00100000;
		color_arr[1372] = 8'b00000000;
		color_arr[1373] = 8'b00000000;
		color_arr[1374] = 8'b00000000;
		color_arr[1375] = 8'b00100000;
		color_arr[1376] = 8'b00100000;
		color_arr[1377] = 8'b00100000;
		color_arr[1378] = 8'b00100000;
		color_arr[1379] = 8'b00100000;
		color_arr[1380] = 8'b00100000;
		color_arr[1381] = 8'b00100000;
		color_arr[1382] = 8'b00100000;
		color_arr[1383] = 8'b00100000;
		color_arr[1384] = 8'b00100000;
		color_arr[1385] = 8'b00100000;
		color_arr[1386] = 8'b00100000;
		color_arr[1387] = 8'b00100000;
		color_arr[1388] = 8'b00000000;
		color_arr[1389] = 8'b00000000;
		color_arr[1390] = 8'b00000000;
		color_arr[1391] = 8'b00000000;
		color_arr[1392] = 8'b00100000;
		color_arr[1393] = 8'b00100000;
		color_arr[1394] = 8'b00100000;
		color_arr[1395] = 8'b00100000;
		color_arr[1396] = 8'b00100000;
		color_arr[1397] = 8'b00100000;
		color_arr[1398] = 8'b00100000;
		color_arr[1399] = 8'b00100000;
		color_arr[1400] = 8'b00100000;
		color_arr[1401] = 8'b00100000;
		color_arr[1402] = 8'b00100000;
		color_arr[1403] = 8'b00100000;
		color_arr[1404] = 8'b00100000;
		color_arr[1405] = 8'b00010010;
		color_arr[1406] = 8'b00010010;
		color_arr[1407] = 8'b00010010;
		color_arr[1408] = 8'b00010010;
		color_arr[1409] = 8'b00010010;
		color_arr[1410] = 8'b00010010;
		color_arr[1411] = 8'b00010010;
		color_arr[1412] = 8'b00010010;
		color_arr[1413] = 8'b00010010;
		color_arr[1414] = 8'b00010010;
		color_arr[1415] = 8'b00010010;
		color_arr[1416] = 8'b00000010;
		color_arr[1417] = 8'b00000010;
		color_arr[1418] = 8'b00000010;
		color_arr[1419] = 8'b00000010;
		color_arr[1420] = 8'b00000010;
		color_arr[1421] = 8'b00000010;
		color_arr[1422] = 8'b00000010;
		color_arr[1423] = 8'b00000010;
		color_arr[1424] = 8'b00000010;
		color_arr[1425] = 8'b00000010;
		color_arr[1426] = 8'b00000010;
		color_arr[1427] = 8'b00000010;
		color_arr[1428] = 8'b00000010;
		color_arr[1429] = 8'b00000010;
		color_arr[1430] = 8'b00000010;
		color_arr[1431] = 8'b00000010;
		color_arr[1432] = 8'b00000010;
		color_arr[1433] = 8'b00000010;
		color_arr[1434] = 8'b00000010;
		color_arr[1435] = 8'b00000010;
		color_arr[1436] = 8'b00000010;
		color_arr[1437] = 8'b00000010;
		color_arr[1438] = 8'b00000010;
		color_arr[1439] = 8'b00000010;
		color_arr[1440] = 8'b00000010;
		color_arr[1441] = 8'b00000010;
		color_arr[1442] = 8'b00000010;
		color_arr[1443] = 8'b00000010;
		color_arr[1444] = 8'b00000010;
		color_arr[1445] = 8'b00000010;
		color_arr[1446] = 8'b00010010;
		color_arr[1447] = 8'b00010010;
		color_arr[1448] = 8'b00000000;
		color_arr[1449] = 8'b00000000;
		color_arr[1450] = 8'b00000000;
		color_arr[1451] = 8'b00000000;
		color_arr[1452] = 8'b00010010;
		color_arr[1453] = 8'b00010010;
		color_arr[1454] = 8'b00010010;
		color_arr[1455] = 8'b00010010;
		color_arr[1456] = 8'b00010010;
		color_arr[1457] = 8'b00010010;
		color_arr[1458] = 8'b00010010;
		color_arr[1459] = 8'b00010010;
		color_arr[1460] = 8'b00010010;
		color_arr[1461] = 8'b00010010;
		color_arr[1462] = 8'b00010010;
		color_arr[1463] = 8'b00010010;
		color_arr[1464] = 8'b00010010;
		color_arr[1465] = 8'b00010010;
		color_arr[1466] = 8'b00010010;
		color_arr[1467] = 8'b00010010;
		color_arr[1468] = 8'b00010010;
		color_arr[1469] = 8'b00010010;
		color_arr[1470] = 8'b00010010;
		color_arr[1471] = 8'b00010010;
		color_arr[1472] = 8'b00010010;
		color_arr[1473] = 8'b00010010;
		color_arr[1474] = 8'b00010010;
		color_arr[1475] = 8'b00010010;
		color_arr[1476] = 8'b00010010;
		color_arr[1477] = 8'b00010010;
		color_arr[1478] = 8'b00010010;
		color_arr[1479] = 8'b00010010;
		color_arr[1480] = 8'b00010010;
		color_arr[1481] = 8'b00010010;
		color_arr[1482] = 8'b00010010;
		color_arr[1483] = 8'b00010010;
		color_arr[1484] = 8'b00010010;
		color_arr[1485] = 8'b00010010;
		color_arr[1486] = 8'b00010010;
		color_arr[1487] = 8'b00010010;
		color_arr[1488] = 8'b00100000;
		color_arr[1489] = 8'b00100000;
		color_arr[1490] = 8'b00100000;
		color_arr[1491] = 8'b00100000;
		color_arr[1492] = 8'b00100000;
		color_arr[1493] = 8'b00100000;
		color_arr[1494] = 8'b00100000;
		color_arr[1495] = 8'b00100000;
		color_arr[1496] = 8'b00100000;
		color_arr[1497] = 8'b00100000;
		color_arr[1498] = 8'b00100000;
		color_arr[1499] = 8'b00100000;
		color_arr[1500] = 8'b00100000;
		color_arr[1501] = 8'b00000000;
		color_arr[1502] = 8'b00000000;
		color_arr[1503] = 8'b00000000;
		color_arr[1504] = 8'b00100000;
		color_arr[1505] = 8'b00100000;
		color_arr[1506] = 8'b00100000;
		color_arr[1507] = 8'b00100000;
		color_arr[1508] = 8'b00100000;
		color_arr[1509] = 8'b00100000;
		color_arr[1510] = 8'b00100000;
		color_arr[1511] = 8'b00100000;
		color_arr[1512] = 8'b00100000;
		color_arr[1513] = 8'b00100000;
		color_arr[1514] = 8'b00100000;
		color_arr[1515] = 8'b00100000;
		color_arr[1516] = 8'b00100000;
		color_arr[1517] = 8'b00000000;
		color_arr[1518] = 8'b00000000;
		color_arr[1519] = 8'b00000000;
		color_arr[1520] = 8'b00000000;
		color_arr[1521] = 8'b00100000;
		color_arr[1522] = 8'b00100000;
		color_arr[1523] = 8'b00100000;
		color_arr[1524] = 8'b00100000;
		color_arr[1525] = 8'b00100000;
		color_arr[1526] = 8'b00100000;
		color_arr[1527] = 8'b00100000;
		color_arr[1528] = 8'b00100000;
		color_arr[1529] = 8'b00100000;
		color_arr[1530] = 8'b00100000;
		color_arr[1531] = 8'b00100000;
		color_arr[1532] = 8'b00100000;
		color_arr[1533] = 8'b00010010;
		color_arr[1534] = 8'b00010010;
		color_arr[1535] = 8'b00010010;
		color_arr[1536] = 8'b00010010;
		color_arr[1537] = 8'b00010010;
		color_arr[1538] = 8'b00010010;
		color_arr[1539] = 8'b00010010;
		color_arr[1540] = 8'b00010010;
		color_arr[1541] = 8'b00010010;
		color_arr[1542] = 8'b00010010;
		color_arr[1543] = 8'b00010010;
		color_arr[1544] = 8'b00000010;
		color_arr[1545] = 8'b00000010;
		color_arr[1546] = 8'b00000010;
		color_arr[1547] = 8'b00000010;
		color_arr[1548] = 8'b00000010;
		color_arr[1549] = 8'b00000010;
		color_arr[1550] = 8'b00000010;
		color_arr[1551] = 8'b00000010;
		color_arr[1552] = 8'b00000010;
		color_arr[1553] = 8'b00000010;
		color_arr[1554] = 8'b00000010;
		color_arr[1555] = 8'b00000010;
		color_arr[1556] = 8'b00000010;
		color_arr[1557] = 8'b00000010;
		color_arr[1558] = 8'b00000010;
		color_arr[1559] = 8'b00000010;
		color_arr[1560] = 8'b00000010;
		color_arr[1561] = 8'b00000010;
		color_arr[1562] = 8'b00000010;
		color_arr[1563] = 8'b00000010;
		color_arr[1564] = 8'b00000010;
		color_arr[1565] = 8'b00000010;
		color_arr[1566] = 8'b00000010;
		color_arr[1567] = 8'b00000010;
		color_arr[1568] = 8'b00000010;
		color_arr[1569] = 8'b00000010;
		color_arr[1570] = 8'b00000010;
		color_arr[1571] = 8'b00000010;
		color_arr[1572] = 8'b00000010;
		color_arr[1573] = 8'b00000010;
		color_arr[1574] = 8'b00010010;
		color_arr[1575] = 8'b00000000;
		color_arr[1576] = 8'b00000000;
		color_arr[1577] = 8'b00000000;
		color_arr[1578] = 8'b00010010;
		color_arr[1579] = 8'b00010010;
		color_arr[1580] = 8'b00010010;
		color_arr[1581] = 8'b00010010;
		color_arr[1582] = 8'b00010010;
		color_arr[1583] = 8'b00010010;
		color_arr[1584] = 8'b00010010;
		color_arr[1585] = 8'b00010010;
		color_arr[1586] = 8'b00010010;
		color_arr[1587] = 8'b00010010;
		color_arr[1588] = 8'b00010010;
		color_arr[1589] = 8'b00010010;
		color_arr[1590] = 8'b00010010;
		color_arr[1591] = 8'b00010010;
		color_arr[1592] = 8'b00010010;
		color_arr[1593] = 8'b00010010;
		color_arr[1594] = 8'b00010010;
		color_arr[1595] = 8'b00010010;
		color_arr[1596] = 8'b00010010;
		color_arr[1597] = 8'b00010010;
		color_arr[1598] = 8'b00010010;
		color_arr[1599] = 8'b00010010;
		color_arr[1600] = 8'b00010010;
		color_arr[1601] = 8'b00010010;
		color_arr[1602] = 8'b00010010;
		color_arr[1603] = 8'b00010010;
		color_arr[1604] = 8'b00010010;
		color_arr[1605] = 8'b00010010;
		color_arr[1606] = 8'b00010010;
		color_arr[1607] = 8'b00010010;
		color_arr[1608] = 8'b00010010;
		color_arr[1609] = 8'b00010010;
		color_arr[1610] = 8'b00010010;
		color_arr[1611] = 8'b00010010;
		color_arr[1612] = 8'b00010010;
		color_arr[1613] = 8'b00010010;
		color_arr[1614] = 8'b00010010;
		color_arr[1615] = 8'b00010010;
		color_arr[1616] = 8'b00100000;
		color_arr[1617] = 8'b00100000;
		color_arr[1618] = 8'b00100000;
		color_arr[1619] = 8'b00100000;
		color_arr[1620] = 8'b00100000;
		color_arr[1621] = 8'b00100000;
		color_arr[1622] = 8'b00100000;
		color_arr[1623] = 8'b00100000;
		color_arr[1624] = 8'b00100000;
		color_arr[1625] = 8'b00100000;
		color_arr[1626] = 8'b00100000;
		color_arr[1627] = 8'b00100000;
		color_arr[1628] = 8'b00100000;
		color_arr[1629] = 8'b00100000;
		color_arr[1630] = 8'b00000000;
		color_arr[1631] = 8'b00000000;
		color_arr[1632] = 8'b00100000;
		color_arr[1633] = 8'b00100000;
		color_arr[1634] = 8'b00100000;
		color_arr[1635] = 8'b00100000;
		color_arr[1636] = 8'b00100000;
		color_arr[1637] = 8'b00100000;
		color_arr[1638] = 8'b00100000;
		color_arr[1639] = 8'b00100000;
		color_arr[1640] = 8'b00100000;
		color_arr[1641] = 8'b00100000;
		color_arr[1642] = 8'b00100000;
		color_arr[1643] = 8'b00100000;
		color_arr[1644] = 8'b00100000;
		color_arr[1645] = 8'b00100000;
		color_arr[1646] = 8'b00100000;
		color_arr[1647] = 8'b00000000;
		color_arr[1648] = 8'b00000000;
		color_arr[1649] = 8'b00000000;
		color_arr[1650] = 8'b00000000;
		color_arr[1651] = 8'b00100000;
		color_arr[1652] = 8'b00100000;
		color_arr[1653] = 8'b00100000;
		color_arr[1654] = 8'b00100000;
		color_arr[1655] = 8'b00100000;
		color_arr[1656] = 8'b00100000;
		color_arr[1657] = 8'b00100000;
		color_arr[1658] = 8'b00100000;
		color_arr[1659] = 8'b00100000;
		color_arr[1660] = 8'b00100000;
		color_arr[1661] = 8'b00010010;
		color_arr[1662] = 8'b00010010;
		color_arr[1663] = 8'b00010010;
		color_arr[1664] = 8'b00010010;
		color_arr[1665] = 8'b00010010;
		color_arr[1666] = 8'b00010010;
		color_arr[1667] = 8'b00010010;
		color_arr[1668] = 8'b00010010;
		color_arr[1669] = 8'b00010010;
		color_arr[1670] = 8'b00010010;
		color_arr[1671] = 8'b00010010;
		color_arr[1672] = 8'b00000010;
		color_arr[1673] = 8'b00000010;
		color_arr[1674] = 8'b00000010;
		color_arr[1675] = 8'b00000010;
		color_arr[1676] = 8'b00000010;
		color_arr[1677] = 8'b00000010;
		color_arr[1678] = 8'b00000010;
		color_arr[1679] = 8'b00000010;
		color_arr[1680] = 8'b00000010;
		color_arr[1681] = 8'b00000010;
		color_arr[1682] = 8'b00000010;
		color_arr[1683] = 8'b00000010;
		color_arr[1684] = 8'b00000010;
		color_arr[1685] = 8'b00000010;
		color_arr[1686] = 8'b00000010;
		color_arr[1687] = 8'b00000010;
		color_arr[1688] = 8'b00000010;
		color_arr[1689] = 8'b00000010;
		color_arr[1690] = 8'b00000010;
		color_arr[1691] = 8'b00000010;
		color_arr[1692] = 8'b00000010;
		color_arr[1693] = 8'b00000010;
		color_arr[1694] = 8'b00000010;
		color_arr[1695] = 8'b00000010;
		color_arr[1696] = 8'b00000010;
		color_arr[1697] = 8'b00000010;
		color_arr[1698] = 8'b00000010;
		color_arr[1699] = 8'b00000010;
		color_arr[1700] = 8'b00000010;
		color_arr[1701] = 8'b00000010;
		color_arr[1702] = 8'b00000000;
		color_arr[1703] = 8'b00000000;
		color_arr[1704] = 8'b00000000;
		color_arr[1705] = 8'b00010010;
		color_arr[1706] = 8'b00010010;
		color_arr[1707] = 8'b00010010;
		color_arr[1708] = 8'b00010010;
		color_arr[1709] = 8'b00010010;
		color_arr[1710] = 8'b00010010;
		color_arr[1711] = 8'b00010010;
		color_arr[1712] = 8'b00010010;
		color_arr[1713] = 8'b00010010;
		color_arr[1714] = 8'b00010010;
		color_arr[1715] = 8'b00010010;
		color_arr[1716] = 8'b00010010;
		color_arr[1717] = 8'b00010010;
		color_arr[1718] = 8'b00010010;
		color_arr[1719] = 8'b00010010;
		color_arr[1720] = 8'b00010010;
		color_arr[1721] = 8'b00010010;
		color_arr[1722] = 8'b00010010;
		color_arr[1723] = 8'b00010010;
		color_arr[1724] = 8'b00010010;
		color_arr[1725] = 8'b00010010;
		color_arr[1726] = 8'b00010010;
		color_arr[1727] = 8'b00010010;
		color_arr[1728] = 8'b00010010;
		color_arr[1729] = 8'b00010010;
		color_arr[1730] = 8'b00010010;
		color_arr[1731] = 8'b00010010;
		color_arr[1732] = 8'b00010010;
		color_arr[1733] = 8'b00010010;
		color_arr[1734] = 8'b00010010;
		color_arr[1735] = 8'b00010010;
		color_arr[1736] = 8'b00010010;
		color_arr[1737] = 8'b00010010;
		color_arr[1738] = 8'b00010010;
		color_arr[1739] = 8'b00010010;
		color_arr[1740] = 8'b00010010;
		color_arr[1741] = 8'b00010010;
		color_arr[1742] = 8'b00010010;
		color_arr[1743] = 8'b00010010;
		color_arr[1744] = 8'b00100000;
		color_arr[1745] = 8'b00100000;
		color_arr[1746] = 8'b00100000;
		color_arr[1747] = 8'b00100000;
		color_arr[1748] = 8'b00100000;
		color_arr[1749] = 8'b00100000;
		color_arr[1750] = 8'b00100000;
		color_arr[1751] = 8'b00100000;
		color_arr[1752] = 8'b00100000;
		color_arr[1753] = 8'b00100000;
		color_arr[1754] = 8'b00100000;
		color_arr[1755] = 8'b00100000;
		color_arr[1756] = 8'b00100000;
		color_arr[1757] = 8'b00100000;
		color_arr[1758] = 8'b00000000;
		color_arr[1759] = 8'b00000000;
		color_arr[1760] = 8'b00000000;
		color_arr[1761] = 8'b00100000;
		color_arr[1762] = 8'b00100000;
		color_arr[1763] = 8'b00100000;
		color_arr[1764] = 8'b00100000;
		color_arr[1765] = 8'b00100000;
		color_arr[1766] = 8'b00100000;
		color_arr[1767] = 8'b00100000;
		color_arr[1768] = 8'b00100000;
		color_arr[1769] = 8'b00100000;
		color_arr[1770] = 8'b00100000;
		color_arr[1771] = 8'b00100000;
		color_arr[1772] = 8'b00100000;
		color_arr[1773] = 8'b00100000;
		color_arr[1774] = 8'b00100000;
		color_arr[1775] = 8'b00100000;
		color_arr[1776] = 8'b00000000;
		color_arr[1777] = 8'b00000000;
		color_arr[1778] = 8'b00000000;
		color_arr[1779] = 8'b00000000;
		color_arr[1780] = 8'b00100000;
		color_arr[1781] = 8'b00100000;
		color_arr[1782] = 8'b00100000;
		color_arr[1783] = 8'b00100000;
		color_arr[1784] = 8'b00100000;
		color_arr[1785] = 8'b00100000;
		color_arr[1786] = 8'b00100000;
		color_arr[1787] = 8'b00100000;
		color_arr[1788] = 8'b00100000;
		color_arr[1789] = 8'b00010010;
		color_arr[1790] = 8'b00010010;
		color_arr[1791] = 8'b00010010;
		color_arr[1792] = 8'b00010010;
		color_arr[1793] = 8'b00010010;
		color_arr[1794] = 8'b00010010;
		color_arr[1795] = 8'b00010010;
		color_arr[1796] = 8'b00010010;
		color_arr[1797] = 8'b00010010;
		color_arr[1798] = 8'b00010010;
		color_arr[1799] = 8'b00010010;
		color_arr[1800] = 8'b00000010;
		color_arr[1801] = 8'b00000010;
		color_arr[1802] = 8'b00000010;
		color_arr[1803] = 8'b00000010;
		color_arr[1804] = 8'b00000010;
		color_arr[1805] = 8'b00000010;
		color_arr[1806] = 8'b00000010;
		color_arr[1807] = 8'b00000010;
		color_arr[1808] = 8'b00000010;
		color_arr[1809] = 8'b00000010;
		color_arr[1810] = 8'b00000010;
		color_arr[1811] = 8'b00000010;
		color_arr[1812] = 8'b00000010;
		color_arr[1813] = 8'b00000010;
		color_arr[1814] = 8'b00000010;
		color_arr[1815] = 8'b00000010;
		color_arr[1816] = 8'b00000010;
		color_arr[1817] = 8'b00000010;
		color_arr[1818] = 8'b00000010;
		color_arr[1819] = 8'b00000010;
		color_arr[1820] = 8'b00000010;
		color_arr[1821] = 8'b00000010;
		color_arr[1822] = 8'b00000010;
		color_arr[1823] = 8'b00000010;
		color_arr[1824] = 8'b00000010;
		color_arr[1825] = 8'b00000010;
		color_arr[1826] = 8'b00000010;
		color_arr[1827] = 8'b00000010;
		color_arr[1828] = 8'b00000000;
		color_arr[1829] = 8'b00000000;
		color_arr[1830] = 8'b00000000;
		color_arr[1831] = 8'b00000000;
		color_arr[1832] = 8'b00010010;
		color_arr[1833] = 8'b00010010;
		color_arr[1834] = 8'b00010010;
		color_arr[1835] = 8'b00010010;
		color_arr[1836] = 8'b00010010;
		color_arr[1837] = 8'b00010010;
		color_arr[1838] = 8'b00010010;
		color_arr[1839] = 8'b00010010;
		color_arr[1840] = 8'b00010010;
		color_arr[1841] = 8'b00010010;
		color_arr[1842] = 8'b00010010;
		color_arr[1843] = 8'b00010010;
		color_arr[1844] = 8'b00010010;
		color_arr[1845] = 8'b00010010;
		color_arr[1846] = 8'b00010010;
		color_arr[1847] = 8'b00010010;
		color_arr[1848] = 8'b00010010;
		color_arr[1849] = 8'b00010010;
		color_arr[1850] = 8'b00010010;
		color_arr[1851] = 8'b00010010;
		color_arr[1852] = 8'b00010010;
		color_arr[1853] = 8'b00010010;
		color_arr[1854] = 8'b00010010;
		color_arr[1855] = 8'b00010010;
		color_arr[1856] = 8'b00010010;
		color_arr[1857] = 8'b00010010;
		color_arr[1858] = 8'b00010010;
		color_arr[1859] = 8'b00010010;
		color_arr[1860] = 8'b00010010;
		color_arr[1861] = 8'b00010010;
		color_arr[1862] = 8'b00010010;
		color_arr[1863] = 8'b00010010;
		color_arr[1864] = 8'b00010010;
		color_arr[1865] = 8'b00010010;
		color_arr[1866] = 8'b00010010;
		color_arr[1867] = 8'b00010010;
		color_arr[1868] = 8'b00010010;
		color_arr[1869] = 8'b00010010;
		color_arr[1870] = 8'b00010010;
		color_arr[1871] = 8'b00010010;
		color_arr[1872] = 8'b00100000;
		color_arr[1873] = 8'b00100000;
		color_arr[1874] = 8'b00100000;
		color_arr[1875] = 8'b00100000;
		color_arr[1876] = 8'b00100000;
		color_arr[1877] = 8'b00100000;
		color_arr[1878] = 8'b00100000;
		color_arr[1879] = 8'b00100000;
		color_arr[1880] = 8'b00100000;
		color_arr[1881] = 8'b00100000;
		color_arr[1882] = 8'b00100000;
		color_arr[1883] = 8'b00100000;
		color_arr[1884] = 8'b00100000;
		color_arr[1885] = 8'b00100000;
		color_arr[1886] = 8'b00100000;
		color_arr[1887] = 8'b00000000;
		color_arr[1888] = 8'b00000000;
		color_arr[1889] = 8'b00100000;
		color_arr[1890] = 8'b00100000;
		color_arr[1891] = 8'b00100000;
		color_arr[1892] = 8'b00100000;
		color_arr[1893] = 8'b00100000;
		color_arr[1894] = 8'b00100000;
		color_arr[1895] = 8'b00100000;
		color_arr[1896] = 8'b00100000;
		color_arr[1897] = 8'b00100000;
		color_arr[1898] = 8'b00100000;
		color_arr[1899] = 8'b00100000;
		color_arr[1900] = 8'b00100000;
		color_arr[1901] = 8'b00100000;
		color_arr[1902] = 8'b00100000;
		color_arr[1903] = 8'b00100000;
		color_arr[1904] = 8'b00100000;
		color_arr[1905] = 8'b00100000;
		color_arr[1906] = 8'b00000000;
		color_arr[1907] = 8'b00000000;
		color_arr[1908] = 8'b00000000;
		color_arr[1909] = 8'b00100000;
		color_arr[1910] = 8'b00100000;
		color_arr[1911] = 8'b00100000;
		color_arr[1912] = 8'b00100000;
		color_arr[1913] = 8'b00100000;
		color_arr[1914] = 8'b00100000;
		color_arr[1915] = 8'b00100000;
		color_arr[1916] = 8'b00100000;
		color_arr[1917] = 8'b00010010;
		color_arr[1918] = 8'b00010010;
		color_arr[1919] = 8'b00010010;
		color_arr[1920] = 8'b00010010;
		color_arr[1921] = 8'b00010010;
		color_arr[1922] = 8'b00010010;
		color_arr[1923] = 8'b00010010;
		color_arr[1924] = 8'b00010010;
		color_arr[1925] = 8'b00010010;
		color_arr[1926] = 8'b00010010;
		color_arr[1927] = 8'b00010010;
		color_arr[1928] = 8'b00000010;
		color_arr[1929] = 8'b00000010;
		color_arr[1930] = 8'b00000010;
		color_arr[1931] = 8'b00000010;
		color_arr[1932] = 8'b00000010;
		color_arr[1933] = 8'b00000010;
		color_arr[1934] = 8'b00000010;
		color_arr[1935] = 8'b00000010;
		color_arr[1936] = 8'b00000010;
		color_arr[1937] = 8'b00000010;
		color_arr[1938] = 8'b00000010;
		color_arr[1939] = 8'b00000010;
		color_arr[1940] = 8'b00000010;
		color_arr[1941] = 8'b00000010;
		color_arr[1942] = 8'b00000010;
		color_arr[1943] = 8'b00000010;
		color_arr[1944] = 8'b00000010;
		color_arr[1945] = 8'b00000010;
		color_arr[1946] = 8'b00000010;
		color_arr[1947] = 8'b00000010;
		color_arr[1948] = 8'b00000010;
		color_arr[1949] = 8'b00000010;
		color_arr[1950] = 8'b00000010;
		color_arr[1951] = 8'b00000010;
		color_arr[1952] = 8'b00000010;
		color_arr[1953] = 8'b00000010;
		color_arr[1954] = 8'b00000010;
		color_arr[1955] = 8'b00000000;
		color_arr[1956] = 8'b00000000;
		color_arr[1957] = 8'b00000000;
		color_arr[1958] = 8'b00000000;
		color_arr[1959] = 8'b00010010;
		color_arr[1960] = 8'b00010010;
		color_arr[1961] = 8'b00010010;
		color_arr[1962] = 8'b00010010;
		color_arr[1963] = 8'b00010010;
		color_arr[1964] = 8'b00010010;
		color_arr[1965] = 8'b00010010;
		color_arr[1966] = 8'b00010010;
		color_arr[1967] = 8'b00010010;
		color_arr[1968] = 8'b00010010;
		color_arr[1969] = 8'b00010010;
		color_arr[1970] = 8'b00010010;
		color_arr[1971] = 8'b00010010;
		color_arr[1972] = 8'b00010010;
		color_arr[1973] = 8'b00010010;
		color_arr[1974] = 8'b00010010;
		color_arr[1975] = 8'b00010010;
		color_arr[1976] = 8'b00010010;
		color_arr[1977] = 8'b00010010;
		color_arr[1978] = 8'b00010010;
		color_arr[1979] = 8'b00010010;
		color_arr[1980] = 8'b00010010;
		color_arr[1981] = 8'b00010010;
		color_arr[1982] = 8'b00010010;
		color_arr[1983] = 8'b00010010;
		color_arr[1984] = 8'b00010010;
		color_arr[1985] = 8'b00010010;
		color_arr[1986] = 8'b00010010;
		color_arr[1987] = 8'b00010010;
		color_arr[1988] = 8'b00010010;
		color_arr[1989] = 8'b00010010;
		color_arr[1990] = 8'b00010010;
		color_arr[1991] = 8'b00010010;
		color_arr[1992] = 8'b00010010;
		color_arr[1993] = 8'b00010010;
		color_arr[1994] = 8'b00010010;
		color_arr[1995] = 8'b00010010;
		color_arr[1996] = 8'b00010010;
		color_arr[1997] = 8'b00010010;
		color_arr[1998] = 8'b00010010;
		color_arr[1999] = 8'b00010010;
		color_arr[2000] = 8'b00100000;
		color_arr[2001] = 8'b00100000;
		color_arr[2002] = 8'b00100000;
		color_arr[2003] = 8'b00100000;
		color_arr[2004] = 8'b00100000;
		color_arr[2005] = 8'b00100000;
		color_arr[2006] = 8'b00100000;
		color_arr[2007] = 8'b00100000;
		color_arr[2008] = 8'b00100000;
		color_arr[2009] = 8'b00100000;
		color_arr[2010] = 8'b00100000;
		color_arr[2011] = 8'b00100000;
		color_arr[2012] = 8'b00100000;
		color_arr[2013] = 8'b00100000;
		color_arr[2014] = 8'b00100000;
		color_arr[2015] = 8'b00000000;
		color_arr[2016] = 8'b00000000;
		color_arr[2017] = 8'b00000000;
		color_arr[2018] = 8'b00100000;
		color_arr[2019] = 8'b00100000;
		color_arr[2020] = 8'b00100000;
		color_arr[2021] = 8'b00100000;
		color_arr[2022] = 8'b00100000;
		color_arr[2023] = 8'b00100000;
		color_arr[2024] = 8'b00100000;
		color_arr[2025] = 8'b00100000;
		color_arr[2026] = 8'b00100000;
		color_arr[2027] = 8'b00100000;
		color_arr[2028] = 8'b00100000;
		color_arr[2029] = 8'b00100000;
		color_arr[2030] = 8'b00100000;
		color_arr[2031] = 8'b00100000;
		color_arr[2032] = 8'b00100000;
		color_arr[2033] = 8'b00100000;
		color_arr[2034] = 8'b00100000;
		color_arr[2035] = 8'b00000000;
		color_arr[2036] = 8'b00000000;
		color_arr[2037] = 8'b00100000;
		color_arr[2038] = 8'b00100000;
		color_arr[2039] = 8'b00100000;
		color_arr[2040] = 8'b00100000;
		color_arr[2041] = 8'b00100000;
		color_arr[2042] = 8'b00100000;
		color_arr[2043] = 8'b00100000;
		color_arr[2044] = 8'b00100000;
		color_arr[2045] = 8'b00010010;
		color_arr[2046] = 8'b00010010;
		color_arr[2047] = 8'b00010010;
		color_arr[2048] = 8'b00010010;
		color_arr[2049] = 8'b00010010;
		color_arr[2050] = 8'b00010010;
		color_arr[2051] = 8'b00010010;
		color_arr[2052] = 8'b00010010;
		color_arr[2053] = 8'b00010010;
		color_arr[2054] = 8'b00010010;
		color_arr[2055] = 8'b00010010;
		color_arr[2056] = 8'b00000010;
		color_arr[2057] = 8'b00000010;
		color_arr[2058] = 8'b00000010;
		color_arr[2059] = 8'b00000010;
		color_arr[2060] = 8'b00000010;
		color_arr[2061] = 8'b00000010;
		color_arr[2062] = 8'b00000010;
		color_arr[2063] = 8'b00000010;
		color_arr[2064] = 8'b00000010;
		color_arr[2065] = 8'b00000010;
		color_arr[2066] = 8'b00000010;
		color_arr[2067] = 8'b00000010;
		color_arr[2068] = 8'b00000010;
		color_arr[2069] = 8'b00000010;
		color_arr[2070] = 8'b00000010;
		color_arr[2071] = 8'b00000010;
		color_arr[2072] = 8'b00000010;
		color_arr[2073] = 8'b00000010;
		color_arr[2074] = 8'b00000010;
		color_arr[2075] = 8'b00000010;
		color_arr[2076] = 8'b00000010;
		color_arr[2077] = 8'b00000010;
		color_arr[2078] = 8'b00000010;
		color_arr[2079] = 8'b00000010;
		color_arr[2080] = 8'b00000010;
		color_arr[2081] = 8'b00000010;
		color_arr[2082] = 8'b00000000;
		color_arr[2083] = 8'b00000000;
		color_arr[2084] = 8'b00000000;
		color_arr[2085] = 8'b00000010;
		color_arr[2086] = 8'b00010010;
		color_arr[2087] = 8'b00010010;
		color_arr[2088] = 8'b00010010;
		color_arr[2089] = 8'b00010010;
		color_arr[2090] = 8'b00010010;
		color_arr[2091] = 8'b00010010;
		color_arr[2092] = 8'b00010010;
		color_arr[2093] = 8'b00010010;
		color_arr[2094] = 8'b00010010;
		color_arr[2095] = 8'b00010010;
		color_arr[2096] = 8'b00010010;
		color_arr[2097] = 8'b00010010;
		color_arr[2098] = 8'b00010010;
		color_arr[2099] = 8'b00010010;
		color_arr[2100] = 8'b00010010;
		color_arr[2101] = 8'b00010010;
		color_arr[2102] = 8'b00010010;
		color_arr[2103] = 8'b00010010;
		color_arr[2104] = 8'b00010010;
		color_arr[2105] = 8'b00010010;
		color_arr[2106] = 8'b00010010;
		color_arr[2107] = 8'b00010010;
		color_arr[2108] = 8'b00010010;
		color_arr[2109] = 8'b00010010;
		color_arr[2110] = 8'b00010010;
		color_arr[2111] = 8'b00010010;
		color_arr[2112] = 8'b00010010;
		color_arr[2113] = 8'b00010010;
		color_arr[2114] = 8'b00010010;
		color_arr[2115] = 8'b00010010;
		color_arr[2116] = 8'b00010010;
		color_arr[2117] = 8'b00010010;
		color_arr[2118] = 8'b00010010;
		color_arr[2119] = 8'b00010010;
		color_arr[2120] = 8'b00010010;
		color_arr[2121] = 8'b00010010;
		color_arr[2122] = 8'b00010010;
		color_arr[2123] = 8'b00010010;
		color_arr[2124] = 8'b00010010;
		color_arr[2125] = 8'b00010010;
		color_arr[2126] = 8'b00010010;
		color_arr[2127] = 8'b00010010;
		color_arr[2128] = 8'b00100000;
		color_arr[2129] = 8'b00100000;
		color_arr[2130] = 8'b00100000;
		color_arr[2131] = 8'b00100000;
		color_arr[2132] = 8'b00100000;
		color_arr[2133] = 8'b00100000;
		color_arr[2134] = 8'b00100000;
		color_arr[2135] = 8'b00100000;
		color_arr[2136] = 8'b00100000;
		color_arr[2137] = 8'b00100000;
		color_arr[2138] = 8'b00100000;
		color_arr[2139] = 8'b00100000;
		color_arr[2140] = 8'b00100000;
		color_arr[2141] = 8'b00100000;
		color_arr[2142] = 8'b00100000;
		color_arr[2143] = 8'b00100000;
		color_arr[2144] = 8'b00000000;
		color_arr[2145] = 8'b00000000;
		color_arr[2146] = 8'b00100000;
		color_arr[2147] = 8'b00100000;
		color_arr[2148] = 8'b00100000;
		color_arr[2149] = 8'b00100000;
		color_arr[2150] = 8'b00100000;
		color_arr[2151] = 8'b00100000;
		color_arr[2152] = 8'b00100000;
		color_arr[2153] = 8'b00100000;
		color_arr[2154] = 8'b00100000;
		color_arr[2155] = 8'b00100000;
		color_arr[2156] = 8'b00100000;
		color_arr[2157] = 8'b00100000;
		color_arr[2158] = 8'b00100000;
		color_arr[2159] = 8'b00100000;
		color_arr[2160] = 8'b00100000;
		color_arr[2161] = 8'b00100000;
		color_arr[2162] = 8'b00100000;
		color_arr[2163] = 8'b00000000;
		color_arr[2164] = 8'b00000000;
		color_arr[2165] = 8'b00000000;
		color_arr[2166] = 8'b00100000;
		color_arr[2167] = 8'b00100000;
		color_arr[2168] = 8'b00100000;
		color_arr[2169] = 8'b00100000;
		color_arr[2170] = 8'b00100000;
		color_arr[2171] = 8'b00100000;
		color_arr[2172] = 8'b00100000;
		color_arr[2173] = 8'b00010010;
		color_arr[2174] = 8'b00010010;
		color_arr[2175] = 8'b00010010;
		color_arr[2176] = 8'b00010010;
		color_arr[2177] = 8'b00010010;
		color_arr[2178] = 8'b00010010;
		color_arr[2179] = 8'b00010010;
		color_arr[2180] = 8'b00010010;
		color_arr[2181] = 8'b00010010;
		color_arr[2182] = 8'b00010010;
		color_arr[2183] = 8'b00010010;
		color_arr[2184] = 8'b00000010;
		color_arr[2185] = 8'b00000010;
		color_arr[2186] = 8'b00000010;
		color_arr[2187] = 8'b00000010;
		color_arr[2188] = 8'b00000010;
		color_arr[2189] = 8'b00000010;
		color_arr[2190] = 8'b00000010;
		color_arr[2191] = 8'b00000010;
		color_arr[2192] = 8'b00000010;
		color_arr[2193] = 8'b00000010;
		color_arr[2194] = 8'b00000010;
		color_arr[2195] = 8'b00000010;
		color_arr[2196] = 8'b00000010;
		color_arr[2197] = 8'b00000010;
		color_arr[2198] = 8'b00000010;
		color_arr[2199] = 8'b00000010;
		color_arr[2200] = 8'b00000010;
		color_arr[2201] = 8'b00000010;
		color_arr[2202] = 8'b00000010;
		color_arr[2203] = 8'b00000010;
		color_arr[2204] = 8'b00000010;
		color_arr[2205] = 8'b00000010;
		color_arr[2206] = 8'b00000010;
		color_arr[2207] = 8'b00000010;
		color_arr[2208] = 8'b00000010;
		color_arr[2209] = 8'b00000000;
		color_arr[2210] = 8'b00000000;
		color_arr[2211] = 8'b00000000;
		color_arr[2212] = 8'b00000010;
		color_arr[2213] = 8'b00000010;
		color_arr[2214] = 8'b00010010;
		color_arr[2215] = 8'b00010010;
		color_arr[2216] = 8'b00010010;
		color_arr[2217] = 8'b00010010;
		color_arr[2218] = 8'b00010010;
		color_arr[2219] = 8'b00010010;
		color_arr[2220] = 8'b00010010;
		color_arr[2221] = 8'b00010010;
		color_arr[2222] = 8'b00010010;
		color_arr[2223] = 8'b00010010;
		color_arr[2224] = 8'b00010010;
		color_arr[2225] = 8'b00010010;
		color_arr[2226] = 8'b00010010;
		color_arr[2227] = 8'b00010010;
		color_arr[2228] = 8'b00010010;
		color_arr[2229] = 8'b00010010;
		color_arr[2230] = 8'b00010010;
		color_arr[2231] = 8'b00010010;
		color_arr[2232] = 8'b00010010;
		color_arr[2233] = 8'b00010010;
		color_arr[2234] = 8'b00010010;
		color_arr[2235] = 8'b00010010;
		color_arr[2236] = 8'b00010010;
		color_arr[2237] = 8'b00010010;
		color_arr[2238] = 8'b00010010;
		color_arr[2239] = 8'b00010010;
		color_arr[2240] = 8'b00010010;
		color_arr[2241] = 8'b00010010;
		color_arr[2242] = 8'b00010010;
		color_arr[2243] = 8'b00010010;
		color_arr[2244] = 8'b00010010;
		color_arr[2245] = 8'b00010010;
		color_arr[2246] = 8'b00010010;
		color_arr[2247] = 8'b00010010;
		color_arr[2248] = 8'b00010010;
		color_arr[2249] = 8'b00010010;
		color_arr[2250] = 8'b00010010;
		color_arr[2251] = 8'b00010010;
		color_arr[2252] = 8'b00010010;
		color_arr[2253] = 8'b00010010;
		color_arr[2254] = 8'b00010010;
		color_arr[2255] = 8'b00010010;
		color_arr[2256] = 8'b00100000;
		color_arr[2257] = 8'b00100000;
		color_arr[2258] = 8'b00100000;
		color_arr[2259] = 8'b00100000;
		color_arr[2260] = 8'b00100000;
		color_arr[2261] = 8'b00100000;
		color_arr[2262] = 8'b00100000;
		color_arr[2263] = 8'b00100000;
		color_arr[2264] = 8'b00100000;
		color_arr[2265] = 8'b00100000;
		color_arr[2266] = 8'b00100000;
		color_arr[2267] = 8'b00100000;
		color_arr[2268] = 8'b00100000;
		color_arr[2269] = 8'b00100000;
		color_arr[2270] = 8'b00100000;
		color_arr[2271] = 8'b00100000;
		color_arr[2272] = 8'b00000000;
		color_arr[2273] = 8'b00000000;
		color_arr[2274] = 8'b00100000;
		color_arr[2275] = 8'b00100000;
		color_arr[2276] = 8'b00100000;
		color_arr[2277] = 8'b00100000;
		color_arr[2278] = 8'b00100000;
		color_arr[2279] = 8'b00100000;
		color_arr[2280] = 8'b00100000;
		color_arr[2281] = 8'b00100000;
		color_arr[2282] = 8'b00100000;
		color_arr[2283] = 8'b00100000;
		color_arr[2284] = 8'b00100000;
		color_arr[2285] = 8'b00100000;
		color_arr[2286] = 8'b00100000;
		color_arr[2287] = 8'b00100000;
		color_arr[2288] = 8'b00100000;
		color_arr[2289] = 8'b00100000;
		color_arr[2290] = 8'b00100000;
		color_arr[2291] = 8'b00100000;
		color_arr[2292] = 8'b00000000;
		color_arr[2293] = 8'b00000000;
		color_arr[2294] = 8'b00000000;
		color_arr[2295] = 8'b00100000;
		color_arr[2296] = 8'b00100000;
		color_arr[2297] = 8'b00100000;
		color_arr[2298] = 8'b00100000;
		color_arr[2299] = 8'b00100000;
		color_arr[2300] = 8'b00100000;
		color_arr[2301] = 8'b00010010;
		color_arr[2302] = 8'b00010010;
		color_arr[2303] = 8'b00010010;
		color_arr[2304] = 8'b00010010;
		color_arr[2305] = 8'b00010010;
		color_arr[2306] = 8'b00010010;
		color_arr[2307] = 8'b00010010;
		color_arr[2308] = 8'b00010010;
		color_arr[2309] = 8'b00010010;
		color_arr[2310] = 8'b00010010;
		color_arr[2311] = 8'b00010010;
		color_arr[2312] = 8'b00000010;
		color_arr[2313] = 8'b00000010;
		color_arr[2314] = 8'b00000010;
		color_arr[2315] = 8'b00000010;
		color_arr[2316] = 8'b00000010;
		color_arr[2317] = 8'b00000010;
		color_arr[2318] = 8'b00000010;
		color_arr[2319] = 8'b00000010;
		color_arr[2320] = 8'b00000010;
		color_arr[2321] = 8'b00000010;
		color_arr[2322] = 8'b00000010;
		color_arr[2323] = 8'b00000010;
		color_arr[2324] = 8'b00000010;
		color_arr[2325] = 8'b00000010;
		color_arr[2326] = 8'b00000010;
		color_arr[2327] = 8'b00000010;
		color_arr[2328] = 8'b00000010;
		color_arr[2329] = 8'b00000010;
		color_arr[2330] = 8'b00000010;
		color_arr[2331] = 8'b00000010;
		color_arr[2332] = 8'b00000010;
		color_arr[2333] = 8'b00000010;
		color_arr[2334] = 8'b00000010;
		color_arr[2335] = 8'b00000010;
		color_arr[2336] = 8'b00000000;
		color_arr[2337] = 8'b00000000;
		color_arr[2338] = 8'b00000000;
		color_arr[2339] = 8'b00000010;
		color_arr[2340] = 8'b00000010;
		color_arr[2341] = 8'b00000010;
		color_arr[2342] = 8'b00010010;
		color_arr[2343] = 8'b00010010;
		color_arr[2344] = 8'b00010010;
		color_arr[2345] = 8'b00010010;
		color_arr[2346] = 8'b00010010;
		color_arr[2347] = 8'b00010010;
		color_arr[2348] = 8'b00010010;
		color_arr[2349] = 8'b00010010;
		color_arr[2350] = 8'b00010010;
		color_arr[2351] = 8'b00010010;
		color_arr[2352] = 8'b00010010;
		color_arr[2353] = 8'b00010010;
		color_arr[2354] = 8'b00010010;
		color_arr[2355] = 8'b00010010;
		color_arr[2356] = 8'b00010010;
		color_arr[2357] = 8'b00010010;
		color_arr[2358] = 8'b00010010;
		color_arr[2359] = 8'b00010010;
		color_arr[2360] = 8'b00010010;
		color_arr[2361] = 8'b00010010;
		color_arr[2362] = 8'b00010010;
		color_arr[2363] = 8'b00010010;
		color_arr[2364] = 8'b00010010;
		color_arr[2365] = 8'b00010010;
		color_arr[2366] = 8'b00010010;
		color_arr[2367] = 8'b00010010;
		color_arr[2368] = 8'b00010010;
		color_arr[2369] = 8'b00010010;
		color_arr[2370] = 8'b00010010;
		color_arr[2371] = 8'b00010010;
		color_arr[2372] = 8'b00010010;
		color_arr[2373] = 8'b00010010;
		color_arr[2374] = 8'b00010010;
		color_arr[2375] = 8'b00010010;
		color_arr[2376] = 8'b00010010;
		color_arr[2377] = 8'b00010010;
		color_arr[2378] = 8'b00010010;
		color_arr[2379] = 8'b00010010;
		color_arr[2380] = 8'b00010010;
		color_arr[2381] = 8'b00010010;
		color_arr[2382] = 8'b00010010;
		color_arr[2383] = 8'b00010010;
		color_arr[2384] = 8'b00100000;
		color_arr[2385] = 8'b00100000;
		color_arr[2386] = 8'b00100000;
		color_arr[2387] = 8'b00100000;
		color_arr[2388] = 8'b00100000;
		color_arr[2389] = 8'b00100000;
		color_arr[2390] = 8'b00100000;
		color_arr[2391] = 8'b00100000;
		color_arr[2392] = 8'b00100000;
		color_arr[2393] = 8'b00100000;
		color_arr[2394] = 8'b00100000;
		color_arr[2395] = 8'b00100000;
		color_arr[2396] = 8'b00100000;
		color_arr[2397] = 8'b00100000;
		color_arr[2398] = 8'b00100000;
		color_arr[2399] = 8'b00100000;
		color_arr[2400] = 8'b00000000;
		color_arr[2401] = 8'b00000000;
		color_arr[2402] = 8'b00000000;
		color_arr[2403] = 8'b00100000;
		color_arr[2404] = 8'b00100000;
		color_arr[2405] = 8'b00100000;
		color_arr[2406] = 8'b00100000;
		color_arr[2407] = 8'b00100000;
		color_arr[2408] = 8'b00100000;
		color_arr[2409] = 8'b00100000;
		color_arr[2410] = 8'b00100000;
		color_arr[2411] = 8'b00100000;
		color_arr[2412] = 8'b00100000;
		color_arr[2413] = 8'b00100000;
		color_arr[2414] = 8'b00100000;
		color_arr[2415] = 8'b00100000;
		color_arr[2416] = 8'b00100000;
		color_arr[2417] = 8'b00100000;
		color_arr[2418] = 8'b00100000;
		color_arr[2419] = 8'b00100000;
		color_arr[2420] = 8'b00100000;
		color_arr[2421] = 8'b00000000;
		color_arr[2422] = 8'b00000000;
		color_arr[2423] = 8'b00100000;
		color_arr[2424] = 8'b00100000;
		color_arr[2425] = 8'b00100000;
		color_arr[2426] = 8'b00100000;
		color_arr[2427] = 8'b00100000;
		color_arr[2428] = 8'b00100000;
		color_arr[2429] = 8'b00010010;
		color_arr[2430] = 8'b00010010;
		color_arr[2431] = 8'b00010010;
		color_arr[2432] = 8'b00010010;
		color_arr[2433] = 8'b00010010;
		color_arr[2434] = 8'b00010010;
		color_arr[2435] = 8'b00010010;
		color_arr[2436] = 8'b00010010;
		color_arr[2437] = 8'b00010010;
		color_arr[2438] = 8'b00010010;
		color_arr[2439] = 8'b00010010;
		color_arr[2440] = 8'b00000010;
		color_arr[2441] = 8'b00000010;
		color_arr[2442] = 8'b00000010;
		color_arr[2443] = 8'b00000010;
		color_arr[2444] = 8'b00000010;
		color_arr[2445] = 8'b00000010;
		color_arr[2446] = 8'b00000010;
		color_arr[2447] = 8'b00000010;
		color_arr[2448] = 8'b00000010;
		color_arr[2449] = 8'b00000010;
		color_arr[2450] = 8'b00000010;
		color_arr[2451] = 8'b00000010;
		color_arr[2452] = 8'b00000010;
		color_arr[2453] = 8'b00000010;
		color_arr[2454] = 8'b00000010;
		color_arr[2455] = 8'b00000010;
		color_arr[2456] = 8'b00000010;
		color_arr[2457] = 8'b00000010;
		color_arr[2458] = 8'b00000010;
		color_arr[2459] = 8'b00000010;
		color_arr[2460] = 8'b00000010;
		color_arr[2461] = 8'b00000010;
		color_arr[2462] = 8'b00000010;
		color_arr[2463] = 8'b00000000;
		color_arr[2464] = 8'b00000000;
		color_arr[2465] = 8'b00000000;
		color_arr[2466] = 8'b00000010;
		color_arr[2467] = 8'b00000010;
		color_arr[2468] = 8'b00000010;
		color_arr[2469] = 8'b00000010;
		color_arr[2470] = 8'b00010010;
		color_arr[2471] = 8'b00010010;
		color_arr[2472] = 8'b00010010;
		color_arr[2473] = 8'b00010010;
		color_arr[2474] = 8'b00010010;
		color_arr[2475] = 8'b00010010;
		color_arr[2476] = 8'b00010010;
		color_arr[2477] = 8'b00010010;
		color_arr[2478] = 8'b00010010;
		color_arr[2479] = 8'b00010010;
		color_arr[2480] = 8'b00010010;
		color_arr[2481] = 8'b00010010;
		color_arr[2482] = 8'b00010010;
		color_arr[2483] = 8'b00010010;
		color_arr[2484] = 8'b00010010;
		color_arr[2485] = 8'b00010010;
		color_arr[2486] = 8'b00010010;
		color_arr[2487] = 8'b00010010;
		color_arr[2488] = 8'b00010010;
		color_arr[2489] = 8'b00010010;
		color_arr[2490] = 8'b00010010;
		color_arr[2491] = 8'b00010010;
		color_arr[2492] = 8'b00010010;
		color_arr[2493] = 8'b00010010;
		color_arr[2494] = 8'b00010010;
		color_arr[2495] = 8'b00010010;
		color_arr[2496] = 8'b00010010;
		color_arr[2497] = 8'b00010010;
		color_arr[2498] = 8'b00010010;
		color_arr[2499] = 8'b00010010;
		color_arr[2500] = 8'b00010010;
		color_arr[2501] = 8'b00010010;
		color_arr[2502] = 8'b00010010;
		color_arr[2503] = 8'b00010010;
		color_arr[2504] = 8'b00010010;
		color_arr[2505] = 8'b00010010;
		color_arr[2506] = 8'b00010010;
		color_arr[2507] = 8'b00010010;
		color_arr[2508] = 8'b00010010;
		color_arr[2509] = 8'b00010010;
		color_arr[2510] = 8'b00010010;
		color_arr[2511] = 8'b00010010;
		color_arr[2512] = 8'b00100000;
		color_arr[2513] = 8'b00100000;
		color_arr[2514] = 8'b00100000;
		color_arr[2515] = 8'b00100000;
		color_arr[2516] = 8'b00100000;
		color_arr[2517] = 8'b00100000;
		color_arr[2518] = 8'b00100000;
		color_arr[2519] = 8'b00100000;
		color_arr[2520] = 8'b00100000;
		color_arr[2521] = 8'b00100000;
		color_arr[2522] = 8'b00100000;
		color_arr[2523] = 8'b00100000;
		color_arr[2524] = 8'b00100000;
		color_arr[2525] = 8'b00100000;
		color_arr[2526] = 8'b00100000;
		color_arr[2527] = 8'b00100000;
		color_arr[2528] = 8'b00100000;
		color_arr[2529] = 8'b00000000;
		color_arr[2530] = 8'b00000000;
		color_arr[2531] = 8'b00100000;
		color_arr[2532] = 8'b00100000;
		color_arr[2533] = 8'b00100000;
		color_arr[2534] = 8'b00100000;
		color_arr[2535] = 8'b00100000;
		color_arr[2536] = 8'b00100000;
		color_arr[2537] = 8'b00100000;
		color_arr[2538] = 8'b00100000;
		color_arr[2539] = 8'b00100000;
		color_arr[2540] = 8'b00100000;
		color_arr[2541] = 8'b00100000;
		color_arr[2542] = 8'b00100000;
		color_arr[2543] = 8'b00100000;
		color_arr[2544] = 8'b00100000;
		color_arr[2545] = 8'b00100000;
		color_arr[2546] = 8'b00100000;
		color_arr[2547] = 8'b00100000;
		color_arr[2548] = 8'b00100000;
		color_arr[2549] = 8'b00000000;
		color_arr[2550] = 8'b00000000;
		color_arr[2551] = 8'b00000000;
		color_arr[2552] = 8'b00100000;
		color_arr[2553] = 8'b00100000;
		color_arr[2554] = 8'b00100000;
		color_arr[2555] = 8'b00100000;
		color_arr[2556] = 8'b00100000;
		color_arr[2557] = 8'b00010010;
		color_arr[2558] = 8'b00010010;
		color_arr[2559] = 8'b00010010;
		color_arr[2560] = 8'b00010010;
		color_arr[2561] = 8'b00010010;
		color_arr[2562] = 8'b00010010;
		color_arr[2563] = 8'b00010010;
		color_arr[2564] = 8'b00010010;
		color_arr[2565] = 8'b00010010;
		color_arr[2566] = 8'b00010010;
		color_arr[2567] = 8'b00010010;
		color_arr[2568] = 8'b00000010;
		color_arr[2569] = 8'b00000010;
		color_arr[2570] = 8'b00000010;
		color_arr[2571] = 8'b00000010;
		color_arr[2572] = 8'b00000010;
		color_arr[2573] = 8'b00000010;
		color_arr[2574] = 8'b00000010;
		color_arr[2575] = 8'b00000010;
		color_arr[2576] = 8'b00000010;
		color_arr[2577] = 8'b00000010;
		color_arr[2578] = 8'b00000010;
		color_arr[2579] = 8'b00000010;
		color_arr[2580] = 8'b00000010;
		color_arr[2581] = 8'b00000010;
		color_arr[2582] = 8'b00000010;
		color_arr[2583] = 8'b00000010;
		color_arr[2584] = 8'b00000010;
		color_arr[2585] = 8'b00000010;
		color_arr[2586] = 8'b00000010;
		color_arr[2587] = 8'b00000010;
		color_arr[2588] = 8'b00000010;
		color_arr[2589] = 8'b00000010;
		color_arr[2590] = 8'b00000000;
		color_arr[2591] = 8'b00000000;
		color_arr[2592] = 8'b00000000;
		color_arr[2593] = 8'b00000010;
		color_arr[2594] = 8'b00000010;
		color_arr[2595] = 8'b00000010;
		color_arr[2596] = 8'b00000010;
		color_arr[2597] = 8'b00000010;
		color_arr[2598] = 8'b00010010;
		color_arr[2599] = 8'b00010010;
		color_arr[2600] = 8'b00010010;
		color_arr[2601] = 8'b00010010;
		color_arr[2602] = 8'b00010010;
		color_arr[2603] = 8'b00010010;
		color_arr[2604] = 8'b00010010;
		color_arr[2605] = 8'b00010010;
		color_arr[2606] = 8'b00010010;
		color_arr[2607] = 8'b00010010;
		color_arr[2608] = 8'b00010010;
		color_arr[2609] = 8'b00010010;
		color_arr[2610] = 8'b00010010;
		color_arr[2611] = 8'b00010010;
		color_arr[2612] = 8'b00010010;
		color_arr[2613] = 8'b00010010;
		color_arr[2614] = 8'b00010010;
		color_arr[2615] = 8'b00010010;
		color_arr[2616] = 8'b00010010;
		color_arr[2617] = 8'b00010010;
		color_arr[2618] = 8'b00010010;
		color_arr[2619] = 8'b00010010;
		color_arr[2620] = 8'b00010010;
		color_arr[2621] = 8'b00010010;
		color_arr[2622] = 8'b00010010;
		color_arr[2623] = 8'b00010010;
		color_arr[2624] = 8'b00010010;
		color_arr[2625] = 8'b00010010;
		color_arr[2626] = 8'b00010010;
		color_arr[2627] = 8'b00010010;
		color_arr[2628] = 8'b00010010;
		color_arr[2629] = 8'b00010010;
		color_arr[2630] = 8'b00010010;
		color_arr[2631] = 8'b00010010;
		color_arr[2632] = 8'b00010010;
		color_arr[2633] = 8'b00010010;
		color_arr[2634] = 8'b00010010;
		color_arr[2635] = 8'b00010010;
		color_arr[2636] = 8'b00010010;
		color_arr[2637] = 8'b00010010;
		color_arr[2638] = 8'b00010010;
		color_arr[2639] = 8'b00010010;
		color_arr[2640] = 8'b00100000;
		color_arr[2641] = 8'b00100000;
		color_arr[2642] = 8'b00100000;
		color_arr[2643] = 8'b00100000;
		color_arr[2644] = 8'b00100000;
		color_arr[2645] = 8'b00100000;
		color_arr[2646] = 8'b00100000;
		color_arr[2647] = 8'b00100000;
		color_arr[2648] = 8'b00100000;
		color_arr[2649] = 8'b00100000;
		color_arr[2650] = 8'b00100000;
		color_arr[2651] = 8'b00100000;
		color_arr[2652] = 8'b00100000;
		color_arr[2653] = 8'b00100000;
		color_arr[2654] = 8'b00100000;
		color_arr[2655] = 8'b00100000;
		color_arr[2656] = 8'b00100000;
		color_arr[2657] = 8'b00000000;
		color_arr[2658] = 8'b00000000;
		color_arr[2659] = 8'b00100000;
		color_arr[2660] = 8'b00100000;
		color_arr[2661] = 8'b00100000;
		color_arr[2662] = 8'b00100000;
		color_arr[2663] = 8'b00100000;
		color_arr[2664] = 8'b00100000;
		color_arr[2665] = 8'b00100000;
		color_arr[2666] = 8'b00100000;
		color_arr[2667] = 8'b00100000;
		color_arr[2668] = 8'b00100000;
		color_arr[2669] = 8'b00100000;
		color_arr[2670] = 8'b00100000;
		color_arr[2671] = 8'b00100000;
		color_arr[2672] = 8'b00100000;
		color_arr[2673] = 8'b00100000;
		color_arr[2674] = 8'b00100000;
		color_arr[2675] = 8'b00100000;
		color_arr[2676] = 8'b00100000;
		color_arr[2677] = 8'b00100000;
		color_arr[2678] = 8'b00000000;
		color_arr[2679] = 8'b00000000;
		color_arr[2680] = 8'b00100000;
		color_arr[2681] = 8'b00100000;
		color_arr[2682] = 8'b00100000;
		color_arr[2683] = 8'b00100000;
		color_arr[2684] = 8'b00100000;
		color_arr[2685] = 8'b00010010;
		color_arr[2686] = 8'b00010010;
		color_arr[2687] = 8'b00010010;
		color_arr[2688] = 8'b00010010;
		color_arr[2689] = 8'b00010010;
		color_arr[2690] = 8'b00010010;
		color_arr[2691] = 8'b00010010;
		color_arr[2692] = 8'b00010010;
		color_arr[2693] = 8'b00010010;
		color_arr[2694] = 8'b00010010;
		color_arr[2695] = 8'b00010010;
		color_arr[2696] = 8'b00000010;
		color_arr[2697] = 8'b00000010;
		color_arr[2698] = 8'b00000010;
		color_arr[2699] = 8'b00000010;
		color_arr[2700] = 8'b00000010;
		color_arr[2701] = 8'b00000010;
		color_arr[2702] = 8'b00000010;
		color_arr[2703] = 8'b00000010;
		color_arr[2704] = 8'b00000010;
		color_arr[2705] = 8'b00000010;
		color_arr[2706] = 8'b00000010;
		color_arr[2707] = 8'b00000010;
		color_arr[2708] = 8'b00000010;
		color_arr[2709] = 8'b00000010;
		color_arr[2710] = 8'b00000010;
		color_arr[2711] = 8'b00000010;
		color_arr[2712] = 8'b00000010;
		color_arr[2713] = 8'b00000010;
		color_arr[2714] = 8'b00000010;
		color_arr[2715] = 8'b00000010;
		color_arr[2716] = 8'b00000010;
		color_arr[2717] = 8'b00000000;
		color_arr[2718] = 8'b00000000;
		color_arr[2719] = 8'b00000000;
		color_arr[2720] = 8'b00000010;
		color_arr[2721] = 8'b00000010;
		color_arr[2722] = 8'b00000010;
		color_arr[2723] = 8'b00000010;
		color_arr[2724] = 8'b00000010;
		color_arr[2725] = 8'b00000010;
		color_arr[2726] = 8'b00010010;
		color_arr[2727] = 8'b00010010;
		color_arr[2728] = 8'b00010010;
		color_arr[2729] = 8'b00010010;
		color_arr[2730] = 8'b00010010;
		color_arr[2731] = 8'b00010010;
		color_arr[2732] = 8'b00010010;
		color_arr[2733] = 8'b00010010;
		color_arr[2734] = 8'b00010010;
		color_arr[2735] = 8'b00010010;
		color_arr[2736] = 8'b00010010;
		color_arr[2737] = 8'b00010010;
		color_arr[2738] = 8'b00010010;
		color_arr[2739] = 8'b00010010;
		color_arr[2740] = 8'b00010010;
		color_arr[2741] = 8'b00010010;
		color_arr[2742] = 8'b00010010;
		color_arr[2743] = 8'b00010010;
		color_arr[2744] = 8'b00010010;
		color_arr[2745] = 8'b00010010;
		color_arr[2746] = 8'b00010010;
		color_arr[2747] = 8'b00010010;
		color_arr[2748] = 8'b00010010;
		color_arr[2749] = 8'b00010010;
		color_arr[2750] = 8'b00010010;
		color_arr[2751] = 8'b00010010;
		color_arr[2752] = 8'b00010010;
		color_arr[2753] = 8'b00010010;
		color_arr[2754] = 8'b00010010;
		color_arr[2755] = 8'b00010010;
		color_arr[2756] = 8'b00010010;
		color_arr[2757] = 8'b00010010;
		color_arr[2758] = 8'b00010010;
		color_arr[2759] = 8'b00010010;
		color_arr[2760] = 8'b00010010;
		color_arr[2761] = 8'b00010010;
		color_arr[2762] = 8'b00010010;
		color_arr[2763] = 8'b00010010;
		color_arr[2764] = 8'b00010010;
		color_arr[2765] = 8'b00010010;
		color_arr[2766] = 8'b00010010;
		color_arr[2767] = 8'b00010010;
		color_arr[2768] = 8'b00100000;
		color_arr[2769] = 8'b00100000;
		color_arr[2770] = 8'b00100000;
		color_arr[2771] = 8'b00100000;
		color_arr[2772] = 8'b00100000;
		color_arr[2773] = 8'b00100000;
		color_arr[2774] = 8'b00100000;
		color_arr[2775] = 8'b00100000;
		color_arr[2776] = 8'b00100000;
		color_arr[2777] = 8'b00100000;
		color_arr[2778] = 8'b00100000;
		color_arr[2779] = 8'b00100000;
		color_arr[2780] = 8'b00100000;
		color_arr[2781] = 8'b00100000;
		color_arr[2782] = 8'b00100000;
		color_arr[2783] = 8'b00100000;
		color_arr[2784] = 8'b00100000;
		color_arr[2785] = 8'b00000000;
		color_arr[2786] = 8'b00000000;
		color_arr[2787] = 8'b00000000;
		color_arr[2788] = 8'b00100000;
		color_arr[2789] = 8'b00100000;
		color_arr[2790] = 8'b00100000;
		color_arr[2791] = 8'b00100000;
		color_arr[2792] = 8'b00100000;
		color_arr[2793] = 8'b00100000;
		color_arr[2794] = 8'b00100000;
		color_arr[2795] = 8'b00100000;
		color_arr[2796] = 8'b00100000;
		color_arr[2797] = 8'b00100000;
		color_arr[2798] = 8'b00100000;
		color_arr[2799] = 8'b00100000;
		color_arr[2800] = 8'b00100000;
		color_arr[2801] = 8'b00100000;
		color_arr[2802] = 8'b00100000;
		color_arr[2803] = 8'b00100000;
		color_arr[2804] = 8'b00100000;
		color_arr[2805] = 8'b00100000;
		color_arr[2806] = 8'b00000000;
		color_arr[2807] = 8'b00000000;
		color_arr[2808] = 8'b00100000;
		color_arr[2809] = 8'b00100000;
		color_arr[2810] = 8'b00100000;
		color_arr[2811] = 8'b00100000;
		color_arr[2812] = 8'b00100000;
		color_arr[2813] = 8'b00010010;
		color_arr[2814] = 8'b00010010;
		color_arr[2815] = 8'b00010010;
		color_arr[2816] = 8'b00010010;
		color_arr[2817] = 8'b00010010;
		color_arr[2818] = 8'b00010010;
		color_arr[2819] = 8'b00010010;
		color_arr[2820] = 8'b00010010;
		color_arr[2821] = 8'b00010010;
		color_arr[2822] = 8'b00010010;
		color_arr[2823] = 8'b00010010;
		color_arr[2824] = 8'b00000010;
		color_arr[2825] = 8'b00000010;
		color_arr[2826] = 8'b00000010;
		color_arr[2827] = 8'b00000010;
		color_arr[2828] = 8'b00000010;
		color_arr[2829] = 8'b00000010;
		color_arr[2830] = 8'b00000010;
		color_arr[2831] = 8'b00000010;
		color_arr[2832] = 8'b00000010;
		color_arr[2833] = 8'b00000010;
		color_arr[2834] = 8'b00000010;
		color_arr[2835] = 8'b00000010;
		color_arr[2836] = 8'b00000010;
		color_arr[2837] = 8'b00000010;
		color_arr[2838] = 8'b00000010;
		color_arr[2839] = 8'b00000010;
		color_arr[2840] = 8'b00000010;
		color_arr[2841] = 8'b00000010;
		color_arr[2842] = 8'b00000010;
		color_arr[2843] = 8'b00000010;
		color_arr[2844] = 8'b00000000;
		color_arr[2845] = 8'b00000000;
		color_arr[2846] = 8'b00000000;
		color_arr[2847] = 8'b00000010;
		color_arr[2848] = 8'b00000010;
		color_arr[2849] = 8'b00000010;
		color_arr[2850] = 8'b00000010;
		color_arr[2851] = 8'b00000010;
		color_arr[2852] = 8'b00000010;
		color_arr[2853] = 8'b00000010;
		color_arr[2854] = 8'b00100000;
		color_arr[2855] = 8'b00100000;
		color_arr[2856] = 8'b00100000;
		color_arr[2857] = 8'b00100000;
		color_arr[2858] = 8'b00100000;
		color_arr[2859] = 8'b00100000;
		color_arr[2860] = 8'b00100000;
		color_arr[2861] = 8'b00100000;
		color_arr[2862] = 8'b00100000;
		color_arr[2863] = 8'b00100000;
		color_arr[2864] = 8'b00100000;
		color_arr[2865] = 8'b00100000;
		color_arr[2866] = 8'b00100000;
		color_arr[2867] = 8'b00100000;
		color_arr[2868] = 8'b00100000;
		color_arr[2869] = 8'b00100000;
		color_arr[2870] = 8'b00100000;
		color_arr[2871] = 8'b00100000;
		color_arr[2872] = 8'b00100000;
		color_arr[2873] = 8'b00100000;
		color_arr[2874] = 8'b00100000;
		color_arr[2875] = 8'b00100000;
		color_arr[2876] = 8'b00100000;
		color_arr[2877] = 8'b00100000;
		color_arr[2878] = 8'b00100000;
		color_arr[2879] = 8'b00100000;
		color_arr[2880] = 8'b00100000;
		color_arr[2881] = 8'b00100000;
		color_arr[2882] = 8'b00100000;
		color_arr[2883] = 8'b00100000;
		color_arr[2884] = 8'b00100000;
		color_arr[2885] = 8'b00100000;
		color_arr[2886] = 8'b00100000;
		color_arr[2887] = 8'b00100000;
		color_arr[2888] = 8'b00100000;
		color_arr[2889] = 8'b00100000;
		color_arr[2890] = 8'b00100000;
		color_arr[2891] = 8'b00100000;
		color_arr[2892] = 8'b00100000;
		color_arr[2893] = 8'b00100000;
		color_arr[2894] = 8'b00100000;
		color_arr[2895] = 8'b00100000;
		color_arr[2896] = 8'b00100000;
		color_arr[2897] = 8'b00100000;
		color_arr[2898] = 8'b00100000;
		color_arr[2899] = 8'b00100000;
		color_arr[2900] = 8'b00100000;
		color_arr[2901] = 8'b00100000;
		color_arr[2902] = 8'b00100000;
		color_arr[2903] = 8'b00100000;
		color_arr[2904] = 8'b00100000;
		color_arr[2905] = 8'b00100000;
		color_arr[2906] = 8'b00100000;
		color_arr[2907] = 8'b00100000;
		color_arr[2908] = 8'b00100000;
		color_arr[2909] = 8'b00100000;
		color_arr[2910] = 8'b00100000;
		color_arr[2911] = 8'b00100000;
		color_arr[2912] = 8'b00100000;
		color_arr[2913] = 8'b00100000;
		color_arr[2914] = 8'b00000000;
		color_arr[2915] = 8'b00000000;
		color_arr[2916] = 8'b00100000;
		color_arr[2917] = 8'b00100000;
		color_arr[2918] = 8'b00100000;
		color_arr[2919] = 8'b00100000;
		color_arr[2920] = 8'b00100000;
		color_arr[2921] = 8'b00100000;
		color_arr[2922] = 8'b00100000;
		color_arr[2923] = 8'b00100000;
		color_arr[2924] = 8'b00100000;
		color_arr[2925] = 8'b00100000;
		color_arr[2926] = 8'b00100000;
		color_arr[2927] = 8'b00100000;
		color_arr[2928] = 8'b00100000;
		color_arr[2929] = 8'b00100000;
		color_arr[2930] = 8'b00100000;
		color_arr[2931] = 8'b00100000;
		color_arr[2932] = 8'b00100000;
		color_arr[2933] = 8'b00100000;
		color_arr[2934] = 8'b00000000;
		color_arr[2935] = 8'b00000000;
		color_arr[2936] = 8'b00000000;
		color_arr[2937] = 8'b00100000;
		color_arr[2938] = 8'b00100000;
		color_arr[2939] = 8'b00100000;
		color_arr[2940] = 8'b00100000;
		color_arr[2941] = 8'b00010010;
		color_arr[2942] = 8'b00010010;
		color_arr[2943] = 8'b00010010;
		color_arr[2944] = 8'b00010010;
		color_arr[2945] = 8'b00010010;
		color_arr[2946] = 8'b00010010;
		color_arr[2947] = 8'b00010010;
		color_arr[2948] = 8'b00010010;
		color_arr[2949] = 8'b00010010;
		color_arr[2950] = 8'b00010010;
		color_arr[2951] = 8'b00010010;
		color_arr[2952] = 8'b00000010;
		color_arr[2953] = 8'b00000010;
		color_arr[2954] = 8'b00000010;
		color_arr[2955] = 8'b00000010;
		color_arr[2956] = 8'b00000010;
		color_arr[2957] = 8'b00000010;
		color_arr[2958] = 8'b00000010;
		color_arr[2959] = 8'b00000010;
		color_arr[2960] = 8'b00000010;
		color_arr[2961] = 8'b00000010;
		color_arr[2962] = 8'b00000010;
		color_arr[2963] = 8'b00000010;
		color_arr[2964] = 8'b00000010;
		color_arr[2965] = 8'b00000010;
		color_arr[2966] = 8'b00000010;
		color_arr[2967] = 8'b00000010;
		color_arr[2968] = 8'b00000010;
		color_arr[2969] = 8'b00000010;
		color_arr[2970] = 8'b00000010;
		color_arr[2971] = 8'b00000000;
		color_arr[2972] = 8'b00000000;
		color_arr[2973] = 8'b00000000;
		color_arr[2974] = 8'b00000010;
		color_arr[2975] = 8'b00000010;
		color_arr[2976] = 8'b00000010;
		color_arr[2977] = 8'b00000010;
		color_arr[2978] = 8'b00000010;
		color_arr[2979] = 8'b00000010;
		color_arr[2980] = 8'b00000010;
		color_arr[2981] = 8'b00000010;
		color_arr[2982] = 8'b00100000;
		color_arr[2983] = 8'b00100000;
		color_arr[2984] = 8'b00100000;
		color_arr[2985] = 8'b00100000;
		color_arr[2986] = 8'b00100000;
		color_arr[2987] = 8'b00100000;
		color_arr[2988] = 8'b00100000;
		color_arr[2989] = 8'b00100000;
		color_arr[2990] = 8'b00100000;
		color_arr[2991] = 8'b00100000;
		color_arr[2992] = 8'b00100000;
		color_arr[2993] = 8'b00100000;
		color_arr[2994] = 8'b00100000;
		color_arr[2995] = 8'b00100000;
		color_arr[2996] = 8'b00100000;
		color_arr[2997] = 8'b00100000;
		color_arr[2998] = 8'b00100000;
		color_arr[2999] = 8'b00100000;
		color_arr[3000] = 8'b00100000;
		color_arr[3001] = 8'b00100000;
		color_arr[3002] = 8'b00100000;
		color_arr[3003] = 8'b00100000;
		color_arr[3004] = 8'b00100000;
		color_arr[3005] = 8'b00100000;
		color_arr[3006] = 8'b00100000;
		color_arr[3007] = 8'b00100000;
		color_arr[3008] = 8'b00100000;
		color_arr[3009] = 8'b00100000;
		color_arr[3010] = 8'b00100000;
		color_arr[3011] = 8'b00100000;
		color_arr[3012] = 8'b00100000;
		color_arr[3013] = 8'b00100000;
		color_arr[3014] = 8'b00100000;
		color_arr[3015] = 8'b00100000;
		color_arr[3016] = 8'b00100000;
		color_arr[3017] = 8'b00100000;
		color_arr[3018] = 8'b00100000;
		color_arr[3019] = 8'b00100000;
		color_arr[3020] = 8'b00100000;
		color_arr[3021] = 8'b00100000;
		color_arr[3022] = 8'b00100000;
		color_arr[3023] = 8'b00100000;
		color_arr[3024] = 8'b00001000;
		color_arr[3025] = 8'b00001000;
		color_arr[3026] = 8'b00001000;
		color_arr[3027] = 8'b00001000;
		color_arr[3028] = 8'b00001000;
		color_arr[3029] = 8'b00001000;
		color_arr[3030] = 8'b00001000;
		color_arr[3031] = 8'b00001000;
		color_arr[3032] = 8'b00001000;
		color_arr[3033] = 8'b00001000;
		color_arr[3034] = 8'b00001000;
		color_arr[3035] = 8'b00001000;
		color_arr[3036] = 8'b00001000;
		color_arr[3037] = 8'b00001000;
		color_arr[3038] = 8'b00001000;
		color_arr[3039] = 8'b00001000;
		color_arr[3040] = 8'b00001000;
		color_arr[3041] = 8'b00001000;
		color_arr[3042] = 8'b00000000;
		color_arr[3043] = 8'b00000000;
		color_arr[3044] = 8'b00001000;
		color_arr[3045] = 8'b00001000;
		color_arr[3046] = 8'b00001000;
		color_arr[3047] = 8'b00001000;
		color_arr[3048] = 8'b00001000;
		color_arr[3049] = 8'b00001000;
		color_arr[3050] = 8'b00001000;
		color_arr[3051] = 8'b00001000;
		color_arr[3052] = 8'b00001000;
		color_arr[3053] = 8'b00001000;
		color_arr[3054] = 8'b00001000;
		color_arr[3055] = 8'b00001000;
		color_arr[3056] = 8'b00001000;
		color_arr[3057] = 8'b00001000;
		color_arr[3058] = 8'b00001000;
		color_arr[3059] = 8'b00001000;
		color_arr[3060] = 8'b00001000;
		color_arr[3061] = 8'b00001000;
		color_arr[3062] = 8'b00001000;
		color_arr[3063] = 8'b00000000;
		color_arr[3064] = 8'b00000000;
		color_arr[3065] = 8'b00001000;
		color_arr[3066] = 8'b00001000;
		color_arr[3067] = 8'b00001000;
		color_arr[3068] = 8'b00001000;
		color_arr[3069] = 8'b00010010;
		color_arr[3070] = 8'b00010010;
		color_arr[3071] = 8'b00010010;
		color_arr[3072] = 8'b00010010;
		color_arr[3073] = 8'b00010010;
		color_arr[3074] = 8'b00010010;
		color_arr[3075] = 8'b00010010;
		color_arr[3076] = 8'b00010010;
		color_arr[3077] = 8'b00010010;
		color_arr[3078] = 8'b00010010;
		color_arr[3079] = 8'b00010010;
		color_arr[3080] = 8'b00000010;
		color_arr[3081] = 8'b00000010;
		color_arr[3082] = 8'b00000010;
		color_arr[3083] = 8'b00000010;
		color_arr[3084] = 8'b00000010;
		color_arr[3085] = 8'b00000010;
		color_arr[3086] = 8'b00000010;
		color_arr[3087] = 8'b00000010;
		color_arr[3088] = 8'b00000010;
		color_arr[3089] = 8'b00000010;
		color_arr[3090] = 8'b00000010;
		color_arr[3091] = 8'b00000010;
		color_arr[3092] = 8'b00000010;
		color_arr[3093] = 8'b00000010;
		color_arr[3094] = 8'b00000010;
		color_arr[3095] = 8'b00000010;
		color_arr[3096] = 8'b00000010;
		color_arr[3097] = 8'b00000010;
		color_arr[3098] = 8'b00000000;
		color_arr[3099] = 8'b00000000;
		color_arr[3100] = 8'b00000000;
		color_arr[3101] = 8'b00000010;
		color_arr[3102] = 8'b00000010;
		color_arr[3103] = 8'b00000010;
		color_arr[3104] = 8'b00000010;
		color_arr[3105] = 8'b00000010;
		color_arr[3106] = 8'b00000010;
		color_arr[3107] = 8'b00000010;
		color_arr[3108] = 8'b00000010;
		color_arr[3109] = 8'b00000010;
		color_arr[3110] = 8'b00100000;
		color_arr[3111] = 8'b00100000;
		color_arr[3112] = 8'b00100000;
		color_arr[3113] = 8'b00100000;
		color_arr[3114] = 8'b00100000;
		color_arr[3115] = 8'b00100000;
		color_arr[3116] = 8'b00100000;
		color_arr[3117] = 8'b00100000;
		color_arr[3118] = 8'b00100000;
		color_arr[3119] = 8'b00100000;
		color_arr[3120] = 8'b00100000;
		color_arr[3121] = 8'b00100000;
		color_arr[3122] = 8'b00100000;
		color_arr[3123] = 8'b00100000;
		color_arr[3124] = 8'b00100000;
		color_arr[3125] = 8'b00100000;
		color_arr[3126] = 8'b00100000;
		color_arr[3127] = 8'b00100000;
		color_arr[3128] = 8'b00100000;
		color_arr[3129] = 8'b00100000;
		color_arr[3130] = 8'b00100000;
		color_arr[3131] = 8'b00100000;
		color_arr[3132] = 8'b00100000;
		color_arr[3133] = 8'b00100000;
		color_arr[3134] = 8'b00100000;
		color_arr[3135] = 8'b00100000;
		color_arr[3136] = 8'b00100000;
		color_arr[3137] = 8'b00100000;
		color_arr[3138] = 8'b00100000;
		color_arr[3139] = 8'b00100000;
		color_arr[3140] = 8'b00100000;
		color_arr[3141] = 8'b00100000;
		color_arr[3142] = 8'b00100000;
		color_arr[3143] = 8'b00100000;
		color_arr[3144] = 8'b00100000;
		color_arr[3145] = 8'b00100000;
		color_arr[3146] = 8'b00100000;
		color_arr[3147] = 8'b00100000;
		color_arr[3148] = 8'b00100000;
		color_arr[3149] = 8'b00100000;
		color_arr[3150] = 8'b00100000;
		color_arr[3151] = 8'b00100000;
		color_arr[3152] = 8'b00001000;
		color_arr[3153] = 8'b00001000;
		color_arr[3154] = 8'b00001000;
		color_arr[3155] = 8'b00001000;
		color_arr[3156] = 8'b00001000;
		color_arr[3157] = 8'b00001000;
		color_arr[3158] = 8'b00001000;
		color_arr[3159] = 8'b00001000;
		color_arr[3160] = 8'b00001000;
		color_arr[3161] = 8'b00001000;
		color_arr[3162] = 8'b00001000;
		color_arr[3163] = 8'b00001000;
		color_arr[3164] = 8'b00001000;
		color_arr[3165] = 8'b00001000;
		color_arr[3166] = 8'b00001000;
		color_arr[3167] = 8'b00001000;
		color_arr[3168] = 8'b00001000;
		color_arr[3169] = 8'b00001000;
		color_arr[3170] = 8'b00000000;
		color_arr[3171] = 8'b00000000;
		color_arr[3172] = 8'b00000000;
		color_arr[3173] = 8'b00001000;
		color_arr[3174] = 8'b00001000;
		color_arr[3175] = 8'b00001000;
		color_arr[3176] = 8'b00001000;
		color_arr[3177] = 8'b00001000;
		color_arr[3178] = 8'b00001000;
		color_arr[3179] = 8'b00001000;
		color_arr[3180] = 8'b00001000;
		color_arr[3181] = 8'b00001000;
		color_arr[3182] = 8'b00001000;
		color_arr[3183] = 8'b00001000;
		color_arr[3184] = 8'b00001000;
		color_arr[3185] = 8'b00001000;
		color_arr[3186] = 8'b00001000;
		color_arr[3187] = 8'b00001000;
		color_arr[3188] = 8'b00001000;
		color_arr[3189] = 8'b00001000;
		color_arr[3190] = 8'b00001000;
		color_arr[3191] = 8'b00000000;
		color_arr[3192] = 8'b00000000;
		color_arr[3193] = 8'b00001000;
		color_arr[3194] = 8'b00001000;
		color_arr[3195] = 8'b00001000;
		color_arr[3196] = 8'b00001000;
		color_arr[3197] = 8'b00010010;
		color_arr[3198] = 8'b00010010;
		color_arr[3199] = 8'b00010010;
		color_arr[3200] = 8'b00010010;
		color_arr[3201] = 8'b00010010;
		color_arr[3202] = 8'b00010010;
		color_arr[3203] = 8'b00010010;
		color_arr[3204] = 8'b00010010;
		color_arr[3205] = 8'b00010010;
		color_arr[3206] = 8'b00010010;
		color_arr[3207] = 8'b00010010;
		color_arr[3208] = 8'b00000010;
		color_arr[3209] = 8'b00000010;
		color_arr[3210] = 8'b00000010;
		color_arr[3211] = 8'b00000010;
		color_arr[3212] = 8'b00000010;
		color_arr[3213] = 8'b00000010;
		color_arr[3214] = 8'b00000010;
		color_arr[3215] = 8'b00000010;
		color_arr[3216] = 8'b00000010;
		color_arr[3217] = 8'b00000010;
		color_arr[3218] = 8'b00000010;
		color_arr[3219] = 8'b00000010;
		color_arr[3220] = 8'b00000010;
		color_arr[3221] = 8'b00000010;
		color_arr[3222] = 8'b00000010;
		color_arr[3223] = 8'b00000010;
		color_arr[3224] = 8'b00000010;
		color_arr[3225] = 8'b00000000;
		color_arr[3226] = 8'b00000000;
		color_arr[3227] = 8'b00000000;
		color_arr[3228] = 8'b00000010;
		color_arr[3229] = 8'b00000010;
		color_arr[3230] = 8'b00000010;
		color_arr[3231] = 8'b00000010;
		color_arr[3232] = 8'b00000010;
		color_arr[3233] = 8'b00000010;
		color_arr[3234] = 8'b00000010;
		color_arr[3235] = 8'b00000010;
		color_arr[3236] = 8'b00000010;
		color_arr[3237] = 8'b00000010;
		color_arr[3238] = 8'b00100000;
		color_arr[3239] = 8'b00100000;
		color_arr[3240] = 8'b00100000;
		color_arr[3241] = 8'b00100000;
		color_arr[3242] = 8'b00100000;
		color_arr[3243] = 8'b00100000;
		color_arr[3244] = 8'b00100000;
		color_arr[3245] = 8'b00100000;
		color_arr[3246] = 8'b00100000;
		color_arr[3247] = 8'b00100000;
		color_arr[3248] = 8'b00100000;
		color_arr[3249] = 8'b00100000;
		color_arr[3250] = 8'b00100000;
		color_arr[3251] = 8'b00100000;
		color_arr[3252] = 8'b00100000;
		color_arr[3253] = 8'b00100000;
		color_arr[3254] = 8'b00100000;
		color_arr[3255] = 8'b00100000;
		color_arr[3256] = 8'b00100000;
		color_arr[3257] = 8'b00100000;
		color_arr[3258] = 8'b00100000;
		color_arr[3259] = 8'b00100000;
		color_arr[3260] = 8'b00100000;
		color_arr[3261] = 8'b00100000;
		color_arr[3262] = 8'b00100000;
		color_arr[3263] = 8'b00100000;
		color_arr[3264] = 8'b00100000;
		color_arr[3265] = 8'b00100000;
		color_arr[3266] = 8'b00100000;
		color_arr[3267] = 8'b00100000;
		color_arr[3268] = 8'b00100000;
		color_arr[3269] = 8'b00100000;
		color_arr[3270] = 8'b00100000;
		color_arr[3271] = 8'b00100000;
		color_arr[3272] = 8'b00100000;
		color_arr[3273] = 8'b00100000;
		color_arr[3274] = 8'b00100000;
		color_arr[3275] = 8'b00100000;
		color_arr[3276] = 8'b00100000;
		color_arr[3277] = 8'b00100000;
		color_arr[3278] = 8'b00100000;
		color_arr[3279] = 8'b00100000;
		color_arr[3280] = 8'b00001000;
		color_arr[3281] = 8'b00001000;
		color_arr[3282] = 8'b00001000;
		color_arr[3283] = 8'b00001000;
		color_arr[3284] = 8'b00001000;
		color_arr[3285] = 8'b00001000;
		color_arr[3286] = 8'b00001000;
		color_arr[3287] = 8'b00001000;
		color_arr[3288] = 8'b00001000;
		color_arr[3289] = 8'b00001000;
		color_arr[3290] = 8'b00001000;
		color_arr[3291] = 8'b00001000;
		color_arr[3292] = 8'b00001000;
		color_arr[3293] = 8'b00001000;
		color_arr[3294] = 8'b00001000;
		color_arr[3295] = 8'b00001000;
		color_arr[3296] = 8'b00001000;
		color_arr[3297] = 8'b00001000;
		color_arr[3298] = 8'b00001000;
		color_arr[3299] = 8'b00000000;
		color_arr[3300] = 8'b00000000;
		color_arr[3301] = 8'b00001000;
		color_arr[3302] = 8'b00001000;
		color_arr[3303] = 8'b00001000;
		color_arr[3304] = 8'b00001000;
		color_arr[3305] = 8'b00001000;
		color_arr[3306] = 8'b00001000;
		color_arr[3307] = 8'b00001000;
		color_arr[3308] = 8'b00001000;
		color_arr[3309] = 8'b00001000;
		color_arr[3310] = 8'b00001000;
		color_arr[3311] = 8'b00001000;
		color_arr[3312] = 8'b00001000;
		color_arr[3313] = 8'b00001000;
		color_arr[3314] = 8'b00001000;
		color_arr[3315] = 8'b00001000;
		color_arr[3316] = 8'b00001000;
		color_arr[3317] = 8'b00001000;
		color_arr[3318] = 8'b00001000;
		color_arr[3319] = 8'b00000000;
		color_arr[3320] = 8'b00000000;
		color_arr[3321] = 8'b00001000;
		color_arr[3322] = 8'b00001000;
		color_arr[3323] = 8'b00001000;
		color_arr[3324] = 8'b00001000;
		color_arr[3325] = 8'b00010010;
		color_arr[3326] = 8'b00010010;
		color_arr[3327] = 8'b00010010;
		color_arr[3328] = 8'b00010010;
		color_arr[3329] = 8'b00010010;
		color_arr[3330] = 8'b00010010;
		color_arr[3331] = 8'b00010010;
		color_arr[3332] = 8'b00010010;
		color_arr[3333] = 8'b00010010;
		color_arr[3334] = 8'b00010010;
		color_arr[3335] = 8'b00010010;
		color_arr[3336] = 8'b00000010;
		color_arr[3337] = 8'b00000010;
		color_arr[3338] = 8'b00000010;
		color_arr[3339] = 8'b00000010;
		color_arr[3340] = 8'b00000010;
		color_arr[3341] = 8'b00000010;
		color_arr[3342] = 8'b00000010;
		color_arr[3343] = 8'b00000010;
		color_arr[3344] = 8'b00000010;
		color_arr[3345] = 8'b00000010;
		color_arr[3346] = 8'b00000010;
		color_arr[3347] = 8'b00000010;
		color_arr[3348] = 8'b00000010;
		color_arr[3349] = 8'b00000010;
		color_arr[3350] = 8'b00000010;
		color_arr[3351] = 8'b00000000;
		color_arr[3352] = 8'b00000000;
		color_arr[3353] = 8'b00000000;
		color_arr[3354] = 8'b00000000;
		color_arr[3355] = 8'b00000010;
		color_arr[3356] = 8'b00000010;
		color_arr[3357] = 8'b00000010;
		color_arr[3358] = 8'b00000010;
		color_arr[3359] = 8'b00000010;
		color_arr[3360] = 8'b00000010;
		color_arr[3361] = 8'b00000010;
		color_arr[3362] = 8'b00000010;
		color_arr[3363] = 8'b00000010;
		color_arr[3364] = 8'b00000010;
		color_arr[3365] = 8'b00000010;
		color_arr[3366] = 8'b00100000;
		color_arr[3367] = 8'b00100000;
		color_arr[3368] = 8'b00100000;
		color_arr[3369] = 8'b00100000;
		color_arr[3370] = 8'b00100000;
		color_arr[3371] = 8'b00100000;
		color_arr[3372] = 8'b00100000;
		color_arr[3373] = 8'b00100000;
		color_arr[3374] = 8'b00100000;
		color_arr[3375] = 8'b00100000;
		color_arr[3376] = 8'b00100000;
		color_arr[3377] = 8'b00100000;
		color_arr[3378] = 8'b00100000;
		color_arr[3379] = 8'b00100000;
		color_arr[3380] = 8'b00100000;
		color_arr[3381] = 8'b00100000;
		color_arr[3382] = 8'b00100000;
		color_arr[3383] = 8'b00100000;
		color_arr[3384] = 8'b00100000;
		color_arr[3385] = 8'b00100000;
		color_arr[3386] = 8'b00100000;
		color_arr[3387] = 8'b00100000;
		color_arr[3388] = 8'b00100000;
		color_arr[3389] = 8'b00100000;
		color_arr[3390] = 8'b00100000;
		color_arr[3391] = 8'b00100000;
		color_arr[3392] = 8'b00100000;
		color_arr[3393] = 8'b00100000;
		color_arr[3394] = 8'b00100000;
		color_arr[3395] = 8'b00100000;
		color_arr[3396] = 8'b00100000;
		color_arr[3397] = 8'b00100000;
		color_arr[3398] = 8'b00100000;
		color_arr[3399] = 8'b00100000;
		color_arr[3400] = 8'b00100000;
		color_arr[3401] = 8'b00100000;
		color_arr[3402] = 8'b00100000;
		color_arr[3403] = 8'b00100000;
		color_arr[3404] = 8'b00100000;
		color_arr[3405] = 8'b00100000;
		color_arr[3406] = 8'b00100000;
		color_arr[3407] = 8'b00100000;
		color_arr[3408] = 8'b00001000;
		color_arr[3409] = 8'b00001000;
		color_arr[3410] = 8'b00001000;
		color_arr[3411] = 8'b00001000;
		color_arr[3412] = 8'b00001000;
		color_arr[3413] = 8'b00001000;
		color_arr[3414] = 8'b00001000;
		color_arr[3415] = 8'b00001000;
		color_arr[3416] = 8'b00001000;
		color_arr[3417] = 8'b00001000;
		color_arr[3418] = 8'b00001000;
		color_arr[3419] = 8'b00001000;
		color_arr[3420] = 8'b00001000;
		color_arr[3421] = 8'b00001000;
		color_arr[3422] = 8'b00001000;
		color_arr[3423] = 8'b00001000;
		color_arr[3424] = 8'b00001000;
		color_arr[3425] = 8'b00001000;
		color_arr[3426] = 8'b00001000;
		color_arr[3427] = 8'b00000000;
		color_arr[3428] = 8'b00000000;
		color_arr[3429] = 8'b00001000;
		color_arr[3430] = 8'b00001000;
		color_arr[3431] = 8'b00001000;
		color_arr[3432] = 8'b00001000;
		color_arr[3433] = 8'b00001000;
		color_arr[3434] = 8'b00001000;
		color_arr[3435] = 8'b00001000;
		color_arr[3436] = 8'b00001000;
		color_arr[3437] = 8'b00001000;
		color_arr[3438] = 8'b00001000;
		color_arr[3439] = 8'b00001000;
		color_arr[3440] = 8'b00001000;
		color_arr[3441] = 8'b00001000;
		color_arr[3442] = 8'b00001000;
		color_arr[3443] = 8'b00001000;
		color_arr[3444] = 8'b00001000;
		color_arr[3445] = 8'b00001000;
		color_arr[3446] = 8'b00001000;
		color_arr[3447] = 8'b00000000;
		color_arr[3448] = 8'b00000000;
		color_arr[3449] = 8'b00001000;
		color_arr[3450] = 8'b00001000;
		color_arr[3451] = 8'b00001000;
		color_arr[3452] = 8'b00001000;
		color_arr[3453] = 8'b00010010;
		color_arr[3454] = 8'b00010010;
		color_arr[3455] = 8'b00010010;
		color_arr[3456] = 8'b00010010;
		color_arr[3457] = 8'b00010010;
		color_arr[3458] = 8'b00010010;
		color_arr[3459] = 8'b00010010;
		color_arr[3460] = 8'b00010010;
		color_arr[3461] = 8'b00010010;
		color_arr[3462] = 8'b00010010;
		color_arr[3463] = 8'b00010010;
		color_arr[3464] = 8'b00000010;
		color_arr[3465] = 8'b00000010;
		color_arr[3466] = 8'b00000010;
		color_arr[3467] = 8'b00000010;
		color_arr[3468] = 8'b00000010;
		color_arr[3469] = 8'b00000010;
		color_arr[3470] = 8'b00000010;
		color_arr[3471] = 8'b00000010;
		color_arr[3472] = 8'b00000010;
		color_arr[3473] = 8'b00000000;
		color_arr[3474] = 8'b00000000;
		color_arr[3475] = 8'b00000000;
		color_arr[3476] = 8'b00000000;
		color_arr[3477] = 8'b00000000;
		color_arr[3478] = 8'b00000000;
		color_arr[3479] = 8'b00000000;
		color_arr[3480] = 8'b00000000;
		color_arr[3481] = 8'b00000000;
		color_arr[3482] = 8'b00000010;
		color_arr[3483] = 8'b00000010;
		color_arr[3484] = 8'b00000010;
		color_arr[3485] = 8'b00000010;
		color_arr[3486] = 8'b00000010;
		color_arr[3487] = 8'b00000010;
		color_arr[3488] = 8'b00000010;
		color_arr[3489] = 8'b00000010;
		color_arr[3490] = 8'b00000010;
		color_arr[3491] = 8'b00000010;
		color_arr[3492] = 8'b00000010;
		color_arr[3493] = 8'b00000010;
		color_arr[3494] = 8'b00100000;
		color_arr[3495] = 8'b00100000;
		color_arr[3496] = 8'b00100000;
		color_arr[3497] = 8'b00100000;
		color_arr[3498] = 8'b00100000;
		color_arr[3499] = 8'b00100000;
		color_arr[3500] = 8'b00100000;
		color_arr[3501] = 8'b00100000;
		color_arr[3502] = 8'b00100000;
		color_arr[3503] = 8'b00100000;
		color_arr[3504] = 8'b00100000;
		color_arr[3505] = 8'b00100000;
		color_arr[3506] = 8'b00100000;
		color_arr[3507] = 8'b00100000;
		color_arr[3508] = 8'b00100000;
		color_arr[3509] = 8'b00100000;
		color_arr[3510] = 8'b00100000;
		color_arr[3511] = 8'b00100000;
		color_arr[3512] = 8'b00100000;
		color_arr[3513] = 8'b00100000;
		color_arr[3514] = 8'b00100000;
		color_arr[3515] = 8'b00100000;
		color_arr[3516] = 8'b00100000;
		color_arr[3517] = 8'b00100000;
		color_arr[3518] = 8'b00100000;
		color_arr[3519] = 8'b00100000;
		color_arr[3520] = 8'b00100000;
		color_arr[3521] = 8'b00100000;
		color_arr[3522] = 8'b00100000;
		color_arr[3523] = 8'b00100000;
		color_arr[3524] = 8'b00100000;
		color_arr[3525] = 8'b00100000;
		color_arr[3526] = 8'b00100000;
		color_arr[3527] = 8'b00100000;
		color_arr[3528] = 8'b00100000;
		color_arr[3529] = 8'b00100000;
		color_arr[3530] = 8'b00100000;
		color_arr[3531] = 8'b00100000;
		color_arr[3532] = 8'b00100000;
		color_arr[3533] = 8'b00100000;
		color_arr[3534] = 8'b00100000;
		color_arr[3535] = 8'b00100000;
		color_arr[3536] = 8'b00001000;
		color_arr[3537] = 8'b00001000;
		color_arr[3538] = 8'b00001000;
		color_arr[3539] = 8'b00001000;
		color_arr[3540] = 8'b00001000;
		color_arr[3541] = 8'b00001000;
		color_arr[3542] = 8'b00001000;
		color_arr[3543] = 8'b00001000;
		color_arr[3544] = 8'b00001000;
		color_arr[3545] = 8'b00001000;
		color_arr[3546] = 8'b00001000;
		color_arr[3547] = 8'b00001000;
		color_arr[3548] = 8'b00001000;
		color_arr[3549] = 8'b00001000;
		color_arr[3550] = 8'b00001000;
		color_arr[3551] = 8'b00001000;
		color_arr[3552] = 8'b00001000;
		color_arr[3553] = 8'b00001000;
		color_arr[3554] = 8'b00001000;
		color_arr[3555] = 8'b00000000;
		color_arr[3556] = 8'b00000000;
		color_arr[3557] = 8'b00001000;
		color_arr[3558] = 8'b00001000;
		color_arr[3559] = 8'b00001000;
		color_arr[3560] = 8'b00001000;
		color_arr[3561] = 8'b00001000;
		color_arr[3562] = 8'b00001000;
		color_arr[3563] = 8'b00001000;
		color_arr[3564] = 8'b00001000;
		color_arr[3565] = 8'b00001000;
		color_arr[3566] = 8'b00001000;
		color_arr[3567] = 8'b00001000;
		color_arr[3568] = 8'b00001000;
		color_arr[3569] = 8'b00001000;
		color_arr[3570] = 8'b00001000;
		color_arr[3571] = 8'b00001000;
		color_arr[3572] = 8'b00001000;
		color_arr[3573] = 8'b00001000;
		color_arr[3574] = 8'b00001000;
		color_arr[3575] = 8'b00000000;
		color_arr[3576] = 8'b00000000;
		color_arr[3577] = 8'b00000000;
		color_arr[3578] = 8'b00001000;
		color_arr[3579] = 8'b00001000;
		color_arr[3580] = 8'b00001000;
		color_arr[3581] = 8'b00010010;
		color_arr[3582] = 8'b00010010;
		color_arr[3583] = 8'b00010010;
		color_arr[3584] = 8'b00010010;
		color_arr[3585] = 8'b00010010;
		color_arr[3586] = 8'b00010010;
		color_arr[3587] = 8'b00010010;
		color_arr[3588] = 8'b00010010;
		color_arr[3589] = 8'b00010010;
		color_arr[3590] = 8'b00010010;
		color_arr[3591] = 8'b00010010;
		color_arr[3592] = 8'b00000010;
		color_arr[3593] = 8'b00000010;
		color_arr[3594] = 8'b00000010;
		color_arr[3595] = 8'b00000010;
		color_arr[3596] = 8'b00000010;
		color_arr[3597] = 8'b00000010;
		color_arr[3598] = 8'b00000010;
		color_arr[3599] = 8'b00000000;
		color_arr[3600] = 8'b00000000;
		color_arr[3601] = 8'b00000000;
		color_arr[3602] = 8'b00000000;
		color_arr[3603] = 8'b00000000;
		color_arr[3604] = 8'b00000000;
		color_arr[3605] = 8'b00000000;
		color_arr[3606] = 8'b00000000;
		color_arr[3607] = 8'b00000000;
		color_arr[3608] = 8'b00000010;
		color_arr[3609] = 8'b00000010;
		color_arr[3610] = 8'b00000010;
		color_arr[3611] = 8'b00000010;
		color_arr[3612] = 8'b00000010;
		color_arr[3613] = 8'b00000010;
		color_arr[3614] = 8'b00000010;
		color_arr[3615] = 8'b00000010;
		color_arr[3616] = 8'b00000010;
		color_arr[3617] = 8'b00000010;
		color_arr[3618] = 8'b00000010;
		color_arr[3619] = 8'b00000010;
		color_arr[3620] = 8'b00000010;
		color_arr[3621] = 8'b00000010;
		color_arr[3622] = 8'b00100000;
		color_arr[3623] = 8'b00100000;
		color_arr[3624] = 8'b00100000;
		color_arr[3625] = 8'b00100000;
		color_arr[3626] = 8'b00100000;
		color_arr[3627] = 8'b00100000;
		color_arr[3628] = 8'b00100000;
		color_arr[3629] = 8'b00100000;
		color_arr[3630] = 8'b00100000;
		color_arr[3631] = 8'b00100000;
		color_arr[3632] = 8'b00100000;
		color_arr[3633] = 8'b00100000;
		color_arr[3634] = 8'b00100000;
		color_arr[3635] = 8'b00100000;
		color_arr[3636] = 8'b00100000;
		color_arr[3637] = 8'b00100000;
		color_arr[3638] = 8'b00100000;
		color_arr[3639] = 8'b00100000;
		color_arr[3640] = 8'b00100000;
		color_arr[3641] = 8'b00100000;
		color_arr[3642] = 8'b00100000;
		color_arr[3643] = 8'b00100000;
		color_arr[3644] = 8'b00100000;
		color_arr[3645] = 8'b00100000;
		color_arr[3646] = 8'b00100000;
		color_arr[3647] = 8'b00100000;
		color_arr[3648] = 8'b00100000;
		color_arr[3649] = 8'b00100000;
		color_arr[3650] = 8'b00100000;
		color_arr[3651] = 8'b00100000;
		color_arr[3652] = 8'b00100000;
		color_arr[3653] = 8'b00100000;
		color_arr[3654] = 8'b00100000;
		color_arr[3655] = 8'b00100000;
		color_arr[3656] = 8'b00100000;
		color_arr[3657] = 8'b00100000;
		color_arr[3658] = 8'b00100000;
		color_arr[3659] = 8'b00100000;
		color_arr[3660] = 8'b00100000;
		color_arr[3661] = 8'b00100000;
		color_arr[3662] = 8'b00100000;
		color_arr[3663] = 8'b00100000;
		color_arr[3664] = 8'b00001000;
		color_arr[3665] = 8'b00001000;
		color_arr[3666] = 8'b00001000;
		color_arr[3667] = 8'b00001000;
		color_arr[3668] = 8'b00001000;
		color_arr[3669] = 8'b00001000;
		color_arr[3670] = 8'b00001000;
		color_arr[3671] = 8'b00001000;
		color_arr[3672] = 8'b00001000;
		color_arr[3673] = 8'b00001000;
		color_arr[3674] = 8'b00001000;
		color_arr[3675] = 8'b00001000;
		color_arr[3676] = 8'b00001000;
		color_arr[3677] = 8'b00001000;
		color_arr[3678] = 8'b00001000;
		color_arr[3679] = 8'b00001000;
		color_arr[3680] = 8'b00001000;
		color_arr[3681] = 8'b00001000;
		color_arr[3682] = 8'b00001000;
		color_arr[3683] = 8'b00000000;
		color_arr[3684] = 8'b00000000;
		color_arr[3685] = 8'b00001000;
		color_arr[3686] = 8'b00001000;
		color_arr[3687] = 8'b00001000;
		color_arr[3688] = 8'b00001000;
		color_arr[3689] = 8'b00001000;
		color_arr[3690] = 8'b00001000;
		color_arr[3691] = 8'b00001000;
		color_arr[3692] = 8'b00001000;
		color_arr[3693] = 8'b00001000;
		color_arr[3694] = 8'b00001000;
		color_arr[3695] = 8'b00001000;
		color_arr[3696] = 8'b00001000;
		color_arr[3697] = 8'b00001000;
		color_arr[3698] = 8'b00001000;
		color_arr[3699] = 8'b00001000;
		color_arr[3700] = 8'b00001000;
		color_arr[3701] = 8'b00001000;
		color_arr[3702] = 8'b00001000;
		color_arr[3703] = 8'b00001000;
		color_arr[3704] = 8'b00000000;
		color_arr[3705] = 8'b00000000;
		color_arr[3706] = 8'b00001000;
		color_arr[3707] = 8'b00001000;
		color_arr[3708] = 8'b00001000;
		color_arr[3709] = 8'b00010010;
		color_arr[3710] = 8'b00010010;
		color_arr[3711] = 8'b00010010;
		color_arr[3712] = 8'b00010010;
		color_arr[3713] = 8'b00010010;
		color_arr[3714] = 8'b00010010;
		color_arr[3715] = 8'b00010010;
		color_arr[3716] = 8'b00010010;
		color_arr[3717] = 8'b00010010;
		color_arr[3718] = 8'b00010010;
		color_arr[3719] = 8'b00010010;
		color_arr[3720] = 8'b00000010;
		color_arr[3721] = 8'b00000010;
		color_arr[3722] = 8'b00000010;
		color_arr[3723] = 8'b00000010;
		color_arr[3724] = 8'b00000010;
		color_arr[3725] = 8'b00000000;
		color_arr[3726] = 8'b00000000;
		color_arr[3727] = 8'b00000000;
		color_arr[3728] = 8'b00000000;
		color_arr[3729] = 8'b00000000;
		color_arr[3730] = 8'b00000010;
		color_arr[3731] = 8'b00000010;
		color_arr[3732] = 8'b00000010;
		color_arr[3733] = 8'b00000000;
		color_arr[3734] = 8'b00000000;
		color_arr[3735] = 8'b00000010;
		color_arr[3736] = 8'b00000010;
		color_arr[3737] = 8'b00000010;
		color_arr[3738] = 8'b00000010;
		color_arr[3739] = 8'b00000010;
		color_arr[3740] = 8'b00000010;
		color_arr[3741] = 8'b00000010;
		color_arr[3742] = 8'b00000010;
		color_arr[3743] = 8'b00000010;
		color_arr[3744] = 8'b00000010;
		color_arr[3745] = 8'b00000010;
		color_arr[3746] = 8'b00000010;
		color_arr[3747] = 8'b00000010;
		color_arr[3748] = 8'b00000010;
		color_arr[3749] = 8'b00000010;
		color_arr[3750] = 8'b00100000;
		color_arr[3751] = 8'b00100000;
		color_arr[3752] = 8'b00100000;
		color_arr[3753] = 8'b00100000;
		color_arr[3754] = 8'b00100000;
		color_arr[3755] = 8'b00100000;
		color_arr[3756] = 8'b00100000;
		color_arr[3757] = 8'b00100000;
		color_arr[3758] = 8'b00100000;
		color_arr[3759] = 8'b00100000;
		color_arr[3760] = 8'b00100000;
		color_arr[3761] = 8'b00100000;
		color_arr[3762] = 8'b00100000;
		color_arr[3763] = 8'b00100000;
		color_arr[3764] = 8'b00100000;
		color_arr[3765] = 8'b00100000;
		color_arr[3766] = 8'b00100000;
		color_arr[3767] = 8'b00100000;
		color_arr[3768] = 8'b00100000;
		color_arr[3769] = 8'b00100000;
		color_arr[3770] = 8'b00100000;
		color_arr[3771] = 8'b00100000;
		color_arr[3772] = 8'b00100000;
		color_arr[3773] = 8'b00100000;
		color_arr[3774] = 8'b00100000;
		color_arr[3775] = 8'b00100000;
		color_arr[3776] = 8'b00100000;
		color_arr[3777] = 8'b00100000;
		color_arr[3778] = 8'b00100000;
		color_arr[3779] = 8'b00100000;
		color_arr[3780] = 8'b00100000;
		color_arr[3781] = 8'b00100000;
		color_arr[3782] = 8'b00100000;
		color_arr[3783] = 8'b00100000;
		color_arr[3784] = 8'b00100000;
		color_arr[3785] = 8'b00100000;
		color_arr[3786] = 8'b00100000;
		color_arr[3787] = 8'b00100000;
		color_arr[3788] = 8'b00100000;
		color_arr[3789] = 8'b00100000;
		color_arr[3790] = 8'b00100000;
		color_arr[3791] = 8'b00100000;
		color_arr[3792] = 8'b00001000;
		color_arr[3793] = 8'b00001000;
		color_arr[3794] = 8'b00001000;
		color_arr[3795] = 8'b00001000;
		color_arr[3796] = 8'b00001000;
		color_arr[3797] = 8'b00001000;
		color_arr[3798] = 8'b00001000;
		color_arr[3799] = 8'b00001000;
		color_arr[3800] = 8'b00001000;
		color_arr[3801] = 8'b00001000;
		color_arr[3802] = 8'b00001000;
		color_arr[3803] = 8'b00001000;
		color_arr[3804] = 8'b00001000;
		color_arr[3805] = 8'b00001000;
		color_arr[3806] = 8'b00001000;
		color_arr[3807] = 8'b00001000;
		color_arr[3808] = 8'b00001000;
		color_arr[3809] = 8'b00001000;
		color_arr[3810] = 8'b00001000;
		color_arr[3811] = 8'b00000000;
		color_arr[3812] = 8'b00000000;
		color_arr[3813] = 8'b00001000;
		color_arr[3814] = 8'b00001000;
		color_arr[3815] = 8'b00001000;
		color_arr[3816] = 8'b00001000;
		color_arr[3817] = 8'b00001000;
		color_arr[3818] = 8'b00001000;
		color_arr[3819] = 8'b00001000;
		color_arr[3820] = 8'b00001000;
		color_arr[3821] = 8'b00001000;
		color_arr[3822] = 8'b00001000;
		color_arr[3823] = 8'b00001000;
		color_arr[3824] = 8'b00001000;
		color_arr[3825] = 8'b00001000;
		color_arr[3826] = 8'b00001000;
		color_arr[3827] = 8'b00001000;
		color_arr[3828] = 8'b00001000;
		color_arr[3829] = 8'b00001000;
		color_arr[3830] = 8'b00001000;
		color_arr[3831] = 8'b00001000;
		color_arr[3832] = 8'b00000000;
		color_arr[3833] = 8'b00000000;
		color_arr[3834] = 8'b00001000;
		color_arr[3835] = 8'b00001000;
		color_arr[3836] = 8'b00001000;
		color_arr[3837] = 8'b00010010;
		color_arr[3838] = 8'b00010010;
		color_arr[3839] = 8'b00010010;
		color_arr[3840] = 8'b00010010;
		color_arr[3841] = 8'b00010010;
		color_arr[3842] = 8'b00010010;
		color_arr[3843] = 8'b00010010;
		color_arr[3844] = 8'b00010010;
		color_arr[3845] = 8'b00010010;
		color_arr[3846] = 8'b00010010;
		color_arr[3847] = 8'b00010010;
		color_arr[3848] = 8'b00000010;
		color_arr[3849] = 8'b00000010;
		color_arr[3850] = 8'b00000010;
		color_arr[3851] = 8'b00000010;
		color_arr[3852] = 8'b00000000;
		color_arr[3853] = 8'b00000000;
		color_arr[3854] = 8'b00000000;
		color_arr[3855] = 8'b00000000;
		color_arr[3856] = 8'b00000010;
		color_arr[3857] = 8'b00000010;
		color_arr[3858] = 8'b00000010;
		color_arr[3859] = 8'b00000010;
		color_arr[3860] = 8'b00000010;
		color_arr[3861] = 8'b00000010;
		color_arr[3862] = 8'b00000010;
		color_arr[3863] = 8'b00000010;
		color_arr[3864] = 8'b00000010;
		color_arr[3865] = 8'b00000010;
		color_arr[3866] = 8'b00000010;
		color_arr[3867] = 8'b00000010;
		color_arr[3868] = 8'b00000010;
		color_arr[3869] = 8'b00000010;
		color_arr[3870] = 8'b00000010;
		color_arr[3871] = 8'b00000010;
		color_arr[3872] = 8'b00000010;
		color_arr[3873] = 8'b00000010;
		color_arr[3874] = 8'b00000010;
		color_arr[3875] = 8'b00000010;
		color_arr[3876] = 8'b00000010;
		color_arr[3877] = 8'b00000010;
		color_arr[3878] = 8'b00100000;
		color_arr[3879] = 8'b00100000;
		color_arr[3880] = 8'b00100000;
		color_arr[3881] = 8'b00100000;
		color_arr[3882] = 8'b00100000;
		color_arr[3883] = 8'b00100000;
		color_arr[3884] = 8'b00100000;
		color_arr[3885] = 8'b00100000;
		color_arr[3886] = 8'b00100000;
		color_arr[3887] = 8'b00100000;
		color_arr[3888] = 8'b00100000;
		color_arr[3889] = 8'b00100000;
		color_arr[3890] = 8'b00100000;
		color_arr[3891] = 8'b00100000;
		color_arr[3892] = 8'b00100000;
		color_arr[3893] = 8'b00100000;
		color_arr[3894] = 8'b00100000;
		color_arr[3895] = 8'b00100000;
		color_arr[3896] = 8'b00100000;
		color_arr[3897] = 8'b00100000;
		color_arr[3898] = 8'b00100000;
		color_arr[3899] = 8'b00100000;
		color_arr[3900] = 8'b00100000;
		color_arr[3901] = 8'b00100000;
		color_arr[3902] = 8'b00100000;
		color_arr[3903] = 8'b00100000;
		color_arr[3904] = 8'b00100000;
		color_arr[3905] = 8'b00100000;
		color_arr[3906] = 8'b00100000;
		color_arr[3907] = 8'b00100000;
		color_arr[3908] = 8'b00100000;
		color_arr[3909] = 8'b00100000;
		color_arr[3910] = 8'b00100000;
		color_arr[3911] = 8'b00100000;
		color_arr[3912] = 8'b00100000;
		color_arr[3913] = 8'b00100000;
		color_arr[3914] = 8'b00100000;
		color_arr[3915] = 8'b00100000;
		color_arr[3916] = 8'b00100000;
		color_arr[3917] = 8'b00100000;
		color_arr[3918] = 8'b00100000;
		color_arr[3919] = 8'b00100000;
		color_arr[3920] = 8'b00001000;
		color_arr[3921] = 8'b00001000;
		color_arr[3922] = 8'b00001000;
		color_arr[3923] = 8'b00001000;
		color_arr[3924] = 8'b00001000;
		color_arr[3925] = 8'b00001000;
		color_arr[3926] = 8'b00001000;
		color_arr[3927] = 8'b00001000;
		color_arr[3928] = 8'b00001000;
		color_arr[3929] = 8'b00001000;
		color_arr[3930] = 8'b00001000;
		color_arr[3931] = 8'b00001000;
		color_arr[3932] = 8'b00001000;
		color_arr[3933] = 8'b00001000;
		color_arr[3934] = 8'b00001000;
		color_arr[3935] = 8'b00001000;
		color_arr[3936] = 8'b00001000;
		color_arr[3937] = 8'b00001000;
		color_arr[3938] = 8'b00000000;
		color_arr[3939] = 8'b00000000;
		color_arr[3940] = 8'b00000000;
		color_arr[3941] = 8'b00001000;
		color_arr[3942] = 8'b00001000;
		color_arr[3943] = 8'b00001000;
		color_arr[3944] = 8'b00001000;
		color_arr[3945] = 8'b00001000;
		color_arr[3946] = 8'b00001000;
		color_arr[3947] = 8'b00001000;
		color_arr[3948] = 8'b00001000;
		color_arr[3949] = 8'b00001000;
		color_arr[3950] = 8'b00001000;
		color_arr[3951] = 8'b00001000;
		color_arr[3952] = 8'b00001000;
		color_arr[3953] = 8'b00001000;
		color_arr[3954] = 8'b00001000;
		color_arr[3955] = 8'b00001000;
		color_arr[3956] = 8'b00001000;
		color_arr[3957] = 8'b00001000;
		color_arr[3958] = 8'b00001000;
		color_arr[3959] = 8'b00001000;
		color_arr[3960] = 8'b00000000;
		color_arr[3961] = 8'b00000000;
		color_arr[3962] = 8'b00001000;
		color_arr[3963] = 8'b00001000;
		color_arr[3964] = 8'b00001000;
		color_arr[3965] = 8'b00010010;
		color_arr[3966] = 8'b00010010;
		color_arr[3967] = 8'b00010010;
		color_arr[3968] = 8'b00010010;
		color_arr[3969] = 8'b00010010;
		color_arr[3970] = 8'b00010010;
		color_arr[3971] = 8'b00010010;
		color_arr[3972] = 8'b00010010;
		color_arr[3973] = 8'b00010010;
		color_arr[3974] = 8'b00010010;
		color_arr[3975] = 8'b00010010;
		color_arr[3976] = 8'b00000010;
		color_arr[3977] = 8'b00000010;
		color_arr[3978] = 8'b00000000;
		color_arr[3979] = 8'b00000000;
		color_arr[3980] = 8'b00000000;
		color_arr[3981] = 8'b00000000;
		color_arr[3982] = 8'b00000010;
		color_arr[3983] = 8'b00000010;
		color_arr[3984] = 8'b00000010;
		color_arr[3985] = 8'b00000010;
		color_arr[3986] = 8'b00000010;
		color_arr[3987] = 8'b00000010;
		color_arr[3988] = 8'b00000010;
		color_arr[3989] = 8'b00000010;
		color_arr[3990] = 8'b00000010;
		color_arr[3991] = 8'b00000010;
		color_arr[3992] = 8'b00000010;
		color_arr[3993] = 8'b00000010;
		color_arr[3994] = 8'b00000010;
		color_arr[3995] = 8'b00000010;
		color_arr[3996] = 8'b00000010;
		color_arr[3997] = 8'b00000010;
		color_arr[3998] = 8'b00000010;
		color_arr[3999] = 8'b00000010;
		color_arr[4000] = 8'b00000010;
		color_arr[4001] = 8'b00000010;
		color_arr[4002] = 8'b00000010;
		color_arr[4003] = 8'b00000010;
		color_arr[4004] = 8'b00000010;
		color_arr[4005] = 8'b00000010;
		color_arr[4006] = 8'b00100000;
		color_arr[4007] = 8'b00100000;
		color_arr[4008] = 8'b00100000;
		color_arr[4009] = 8'b00100000;
		color_arr[4010] = 8'b00100000;
		color_arr[4011] = 8'b00100000;
		color_arr[4012] = 8'b00100000;
		color_arr[4013] = 8'b00100000;
		color_arr[4014] = 8'b00100000;
		color_arr[4015] = 8'b00100000;
		color_arr[4016] = 8'b00100000;
		color_arr[4017] = 8'b00100000;
		color_arr[4018] = 8'b00100000;
		color_arr[4019] = 8'b00100000;
		color_arr[4020] = 8'b00100000;
		color_arr[4021] = 8'b00100000;
		color_arr[4022] = 8'b00000000;
		color_arr[4023] = 8'b00000000;
		color_arr[4024] = 8'b00000000;
		color_arr[4025] = 8'b00000000;
		color_arr[4026] = 8'b00000000;
		color_arr[4027] = 8'b00000000;
		color_arr[4028] = 8'b00000000;
		color_arr[4029] = 8'b00000000;
		color_arr[4030] = 8'b00000000;
		color_arr[4031] = 8'b00000000;
		color_arr[4032] = 8'b00000000;
		color_arr[4033] = 8'b00100000;
		color_arr[4034] = 8'b00100000;
		color_arr[4035] = 8'b00100000;
		color_arr[4036] = 8'b00100000;
		color_arr[4037] = 8'b00100000;
		color_arr[4038] = 8'b00100000;
		color_arr[4039] = 8'b00100000;
		color_arr[4040] = 8'b00100000;
		color_arr[4041] = 8'b00100000;
		color_arr[4042] = 8'b00100000;
		color_arr[4043] = 8'b00100000;
		color_arr[4044] = 8'b00100000;
		color_arr[4045] = 8'b00100000;
		color_arr[4046] = 8'b00100000;
		color_arr[4047] = 8'b00100000;
		color_arr[4048] = 8'b00001000;
		color_arr[4049] = 8'b00001000;
		color_arr[4050] = 8'b00001000;
		color_arr[4051] = 8'b00001000;
		color_arr[4052] = 8'b00001000;
		color_arr[4053] = 8'b00001000;
		color_arr[4054] = 8'b00001000;
		color_arr[4055] = 8'b00001000;
		color_arr[4056] = 8'b00001000;
		color_arr[4057] = 8'b00001000;
		color_arr[4058] = 8'b00001000;
		color_arr[4059] = 8'b00001000;
		color_arr[4060] = 8'b00001000;
		color_arr[4061] = 8'b00001000;
		color_arr[4062] = 8'b00001000;
		color_arr[4063] = 8'b00001000;
		color_arr[4064] = 8'b00001000;
		color_arr[4065] = 8'b00000000;
		color_arr[4066] = 8'b00000000;
		color_arr[4067] = 8'b00000000;
		color_arr[4068] = 8'b00001000;
		color_arr[4069] = 8'b00001000;
		color_arr[4070] = 8'b00001000;
		color_arr[4071] = 8'b00001000;
		color_arr[4072] = 8'b00001000;
		color_arr[4073] = 8'b00001000;
		color_arr[4074] = 8'b00001000;
		color_arr[4075] = 8'b00001000;
		color_arr[4076] = 8'b00001000;
		color_arr[4077] = 8'b00001000;
		color_arr[4078] = 8'b00001000;
		color_arr[4079] = 8'b00001000;
		color_arr[4080] = 8'b00001000;
		color_arr[4081] = 8'b00001000;
		color_arr[4082] = 8'b00001000;
		color_arr[4083] = 8'b00001000;
		color_arr[4084] = 8'b00001000;
		color_arr[4085] = 8'b00001000;
		color_arr[4086] = 8'b00001000;
		color_arr[4087] = 8'b00001000;
		color_arr[4088] = 8'b00000000;
		color_arr[4089] = 8'b00000000;
		color_arr[4090] = 8'b00001000;
		color_arr[4091] = 8'b00001000;
		color_arr[4092] = 8'b00001000;
		color_arr[4093] = 8'b00010010;
		color_arr[4094] = 8'b00010010;
		color_arr[4095] = 8'b00010010;
		color_arr[4096] = 8'b00010010;
		color_arr[4097] = 8'b00010010;
		color_arr[4098] = 8'b00010010;
		color_arr[4099] = 8'b00010010;
		color_arr[4100] = 8'b00010010;
		color_arr[4101] = 8'b00010010;
		color_arr[4102] = 8'b00010010;
		color_arr[4103] = 8'b00010010;
		color_arr[4104] = 8'b00000010;
		color_arr[4105] = 8'b00000000;
		color_arr[4106] = 8'b00000000;
		color_arr[4107] = 8'b00000000;
		color_arr[4108] = 8'b00000000;
		color_arr[4109] = 8'b00000010;
		color_arr[4110] = 8'b00000010;
		color_arr[4111] = 8'b00000010;
		color_arr[4112] = 8'b00000010;
		color_arr[4113] = 8'b00000010;
		color_arr[4114] = 8'b00000010;
		color_arr[4115] = 8'b00000010;
		color_arr[4116] = 8'b00000010;
		color_arr[4117] = 8'b00000010;
		color_arr[4118] = 8'b00000010;
		color_arr[4119] = 8'b00000010;
		color_arr[4120] = 8'b00000010;
		color_arr[4121] = 8'b00000010;
		color_arr[4122] = 8'b00000010;
		color_arr[4123] = 8'b00000010;
		color_arr[4124] = 8'b00000010;
		color_arr[4125] = 8'b00000010;
		color_arr[4126] = 8'b00000010;
		color_arr[4127] = 8'b00000010;
		color_arr[4128] = 8'b00000010;
		color_arr[4129] = 8'b00000010;
		color_arr[4130] = 8'b00000010;
		color_arr[4131] = 8'b00000010;
		color_arr[4132] = 8'b00000010;
		color_arr[4133] = 8'b00000010;
		color_arr[4134] = 8'b00100000;
		color_arr[4135] = 8'b00100000;
		color_arr[4136] = 8'b00100000;
		color_arr[4137] = 8'b00100000;
		color_arr[4138] = 8'b00100000;
		color_arr[4139] = 8'b00100000;
		color_arr[4140] = 8'b00100000;
		color_arr[4141] = 8'b00100000;
		color_arr[4142] = 8'b00100000;
		color_arr[4143] = 8'b00100000;
		color_arr[4144] = 8'b00000000;
		color_arr[4145] = 8'b00000000;
		color_arr[4146] = 8'b00000000;
		color_arr[4147] = 8'b00000000;
		color_arr[4148] = 8'b00000000;
		color_arr[4149] = 8'b00000000;
		color_arr[4150] = 8'b00000000;
		color_arr[4151] = 8'b00000000;
		color_arr[4152] = 8'b00000000;
		color_arr[4153] = 8'b00000000;
		color_arr[4154] = 8'b00000000;
		color_arr[4155] = 8'b00000000;
		color_arr[4156] = 8'b00000000;
		color_arr[4157] = 8'b00000000;
		color_arr[4158] = 8'b00000000;
		color_arr[4159] = 8'b00000000;
		color_arr[4160] = 8'b00000000;
		color_arr[4161] = 8'b00000000;
		color_arr[4162] = 8'b00000000;
		color_arr[4163] = 8'b00000000;
		color_arr[4164] = 8'b00000000;
		color_arr[4165] = 8'b00000000;
		color_arr[4166] = 8'b00000000;
		color_arr[4167] = 8'b00000000;
		color_arr[4168] = 8'b00000000;
		color_arr[4169] = 8'b00000000;
		color_arr[4170] = 8'b00000000;
		color_arr[4171] = 8'b00100000;
		color_arr[4172] = 8'b00100000;
		color_arr[4173] = 8'b00100000;
		color_arr[4174] = 8'b00100000;
		color_arr[4175] = 8'b00100000;
		color_arr[4176] = 8'b00001000;
		color_arr[4177] = 8'b00001000;
		color_arr[4178] = 8'b00001000;
		color_arr[4179] = 8'b00001000;
		color_arr[4180] = 8'b00001000;
		color_arr[4181] = 8'b00001000;
		color_arr[4182] = 8'b00001000;
		color_arr[4183] = 8'b00001000;
		color_arr[4184] = 8'b00001000;
		color_arr[4185] = 8'b00001000;
		color_arr[4186] = 8'b00001000;
		color_arr[4187] = 8'b00001000;
		color_arr[4188] = 8'b00001000;
		color_arr[4189] = 8'b00001000;
		color_arr[4190] = 8'b00001000;
		color_arr[4191] = 8'b00001000;
		color_arr[4192] = 8'b00000000;
		color_arr[4193] = 8'b00000000;
		color_arr[4194] = 8'b00000000;
		color_arr[4195] = 8'b00001000;
		color_arr[4196] = 8'b00001000;
		color_arr[4197] = 8'b00001000;
		color_arr[4198] = 8'b00001000;
		color_arr[4199] = 8'b00001000;
		color_arr[4200] = 8'b00001000;
		color_arr[4201] = 8'b00001000;
		color_arr[4202] = 8'b00001000;
		color_arr[4203] = 8'b00001000;
		color_arr[4204] = 8'b00001000;
		color_arr[4205] = 8'b00001000;
		color_arr[4206] = 8'b00001000;
		color_arr[4207] = 8'b00001000;
		color_arr[4208] = 8'b00001000;
		color_arr[4209] = 8'b00001000;
		color_arr[4210] = 8'b00001000;
		color_arr[4211] = 8'b00001000;
		color_arr[4212] = 8'b00001000;
		color_arr[4213] = 8'b00001000;
		color_arr[4214] = 8'b00001000;
		color_arr[4215] = 8'b00000000;
		color_arr[4216] = 8'b00000000;
		color_arr[4217] = 8'b00000000;
		color_arr[4218] = 8'b00001000;
		color_arr[4219] = 8'b00001000;
		color_arr[4220] = 8'b00001000;
		color_arr[4221] = 8'b00010010;
		color_arr[4222] = 8'b00010010;
		color_arr[4223] = 8'b00010010;
		color_arr[4224] = 8'b00010010;
		color_arr[4225] = 8'b00010010;
		color_arr[4226] = 8'b00010010;
		color_arr[4227] = 8'b00010010;
		color_arr[4228] = 8'b00010010;
		color_arr[4229] = 8'b00010010;
		color_arr[4230] = 8'b00010010;
		color_arr[4231] = 8'b00010010;
		color_arr[4232] = 8'b00000000;
		color_arr[4233] = 8'b00000000;
		color_arr[4234] = 8'b00000000;
		color_arr[4235] = 8'b00000010;
		color_arr[4236] = 8'b00000010;
		color_arr[4237] = 8'b00000010;
		color_arr[4238] = 8'b00000010;
		color_arr[4239] = 8'b00000010;
		color_arr[4240] = 8'b00000010;
		color_arr[4241] = 8'b00000010;
		color_arr[4242] = 8'b00000010;
		color_arr[4243] = 8'b00000010;
		color_arr[4244] = 8'b00000010;
		color_arr[4245] = 8'b00000010;
		color_arr[4246] = 8'b00000010;
		color_arr[4247] = 8'b00000010;
		color_arr[4248] = 8'b00000010;
		color_arr[4249] = 8'b00000010;
		color_arr[4250] = 8'b00000010;
		color_arr[4251] = 8'b00000010;
		color_arr[4252] = 8'b00000010;
		color_arr[4253] = 8'b00000010;
		color_arr[4254] = 8'b00000010;
		color_arr[4255] = 8'b00000010;
		color_arr[4256] = 8'b00000010;
		color_arr[4257] = 8'b00000010;
		color_arr[4258] = 8'b00000010;
		color_arr[4259] = 8'b00000010;
		color_arr[4260] = 8'b00000010;
		color_arr[4261] = 8'b00000010;
		color_arr[4262] = 8'b00100000;
		color_arr[4263] = 8'b00100000;
		color_arr[4264] = 8'b00100000;
		color_arr[4265] = 8'b00100000;
		color_arr[4266] = 8'b00100000;
		color_arr[4267] = 8'b00000000;
		color_arr[4268] = 8'b00000000;
		color_arr[4269] = 8'b00000000;
		color_arr[4270] = 8'b00000000;
		color_arr[4271] = 8'b00000000;
		color_arr[4272] = 8'b00000000;
		color_arr[4273] = 8'b00000000;
		color_arr[4274] = 8'b00000000;
		color_arr[4275] = 8'b00000000;
		color_arr[4276] = 8'b00000000;
		color_arr[4277] = 8'b00000000;
		color_arr[4278] = 8'b00000000;
		color_arr[4279] = 8'b00100000;
		color_arr[4280] = 8'b00100000;
		color_arr[4281] = 8'b00100000;
		color_arr[4282] = 8'b00100000;
		color_arr[4283] = 8'b00100000;
		color_arr[4284] = 8'b00100000;
		color_arr[4285] = 8'b00100000;
		color_arr[4286] = 8'b00100000;
		color_arr[4287] = 8'b00100000;
		color_arr[4288] = 8'b00000000;
		color_arr[4289] = 8'b00000000;
		color_arr[4290] = 8'b00000000;
		color_arr[4291] = 8'b00000000;
		color_arr[4292] = 8'b00000000;
		color_arr[4293] = 8'b00000000;
		color_arr[4294] = 8'b00000000;
		color_arr[4295] = 8'b00000000;
		color_arr[4296] = 8'b00000000;
		color_arr[4297] = 8'b00000000;
		color_arr[4298] = 8'b00000000;
		color_arr[4299] = 8'b00000000;
		color_arr[4300] = 8'b00000000;
		color_arr[4301] = 8'b00000000;
		color_arr[4302] = 8'b00000000;
		color_arr[4303] = 8'b00000000;
		color_arr[4304] = 8'b00000000;
		color_arr[4305] = 8'b00001000;
		color_arr[4306] = 8'b00001000;
		color_arr[4307] = 8'b00001000;
		color_arr[4308] = 8'b00001000;
		color_arr[4309] = 8'b00001000;
		color_arr[4310] = 8'b00001000;
		color_arr[4311] = 8'b00001000;
		color_arr[4312] = 8'b00001000;
		color_arr[4313] = 8'b00001000;
		color_arr[4314] = 8'b00001000;
		color_arr[4315] = 8'b00001000;
		color_arr[4316] = 8'b00001000;
		color_arr[4317] = 8'b00001000;
		color_arr[4318] = 8'b00001000;
		color_arr[4319] = 8'b00001000;
		color_arr[4320] = 8'b00000000;
		color_arr[4321] = 8'b00000000;
		color_arr[4322] = 8'b00001000;
		color_arr[4323] = 8'b00001000;
		color_arr[4324] = 8'b00001000;
		color_arr[4325] = 8'b00001000;
		color_arr[4326] = 8'b00001000;
		color_arr[4327] = 8'b00001000;
		color_arr[4328] = 8'b00001000;
		color_arr[4329] = 8'b00001000;
		color_arr[4330] = 8'b00001000;
		color_arr[4331] = 8'b00001000;
		color_arr[4332] = 8'b00001000;
		color_arr[4333] = 8'b00001000;
		color_arr[4334] = 8'b00001000;
		color_arr[4335] = 8'b00001000;
		color_arr[4336] = 8'b00001000;
		color_arr[4337] = 8'b00001000;
		color_arr[4338] = 8'b00001000;
		color_arr[4339] = 8'b00001000;
		color_arr[4340] = 8'b00001000;
		color_arr[4341] = 8'b00001000;
		color_arr[4342] = 8'b00001000;
		color_arr[4343] = 8'b00000000;
		color_arr[4344] = 8'b00000000;
		color_arr[4345] = 8'b00001000;
		color_arr[4346] = 8'b00001000;
		color_arr[4347] = 8'b00001000;
		color_arr[4348] = 8'b00001000;
		color_arr[4349] = 8'b00010010;
		color_arr[4350] = 8'b00010010;
		color_arr[4351] = 8'b00010010;
		color_arr[4352] = 8'b00010010;
		color_arr[4353] = 8'b00010010;
		color_arr[4354] = 8'b00010010;
		color_arr[4355] = 8'b00010010;
		color_arr[4356] = 8'b00010010;
		color_arr[4357] = 8'b00010010;
		color_arr[4358] = 8'b00010010;
		color_arr[4359] = 8'b00000000;
		color_arr[4360] = 8'b00000000;
		color_arr[4361] = 8'b00000000;
		color_arr[4362] = 8'b00000010;
		color_arr[4363] = 8'b00000010;
		color_arr[4364] = 8'b00000010;
		color_arr[4365] = 8'b00000010;
		color_arr[4366] = 8'b00000010;
		color_arr[4367] = 8'b00000010;
		color_arr[4368] = 8'b00000010;
		color_arr[4369] = 8'b00000010;
		color_arr[4370] = 8'b00000010;
		color_arr[4371] = 8'b00000010;
		color_arr[4372] = 8'b00000010;
		color_arr[4373] = 8'b00000010;
		color_arr[4374] = 8'b00000010;
		color_arr[4375] = 8'b00000010;
		color_arr[4376] = 8'b00000010;
		color_arr[4377] = 8'b00000010;
		color_arr[4378] = 8'b00000010;
		color_arr[4379] = 8'b00000010;
		color_arr[4380] = 8'b00000010;
		color_arr[4381] = 8'b00000010;
		color_arr[4382] = 8'b00000010;
		color_arr[4383] = 8'b00000010;
		color_arr[4384] = 8'b00000010;
		color_arr[4385] = 8'b00000010;
		color_arr[4386] = 8'b00000010;
		color_arr[4387] = 8'b00000010;
		color_arr[4388] = 8'b00000010;
		color_arr[4389] = 8'b00000010;
		color_arr[4390] = 8'b00100000;
		color_arr[4391] = 8'b00000000;
		color_arr[4392] = 8'b00000000;
		color_arr[4393] = 8'b00000000;
		color_arr[4394] = 8'b00000000;
		color_arr[4395] = 8'b00000000;
		color_arr[4396] = 8'b00000000;
		color_arr[4397] = 8'b00000000;
		color_arr[4398] = 8'b00000000;
		color_arr[4399] = 8'b00000000;
		color_arr[4400] = 8'b00000000;
		color_arr[4401] = 8'b00100000;
		color_arr[4402] = 8'b00100000;
		color_arr[4403] = 8'b00100000;
		color_arr[4404] = 8'b00100000;
		color_arr[4405] = 8'b00100000;
		color_arr[4406] = 8'b00100000;
		color_arr[4407] = 8'b00100000;
		color_arr[4408] = 8'b00100000;
		color_arr[4409] = 8'b00100000;
		color_arr[4410] = 8'b00100000;
		color_arr[4411] = 8'b00100000;
		color_arr[4412] = 8'b00100000;
		color_arr[4413] = 8'b00100000;
		color_arr[4414] = 8'b00100000;
		color_arr[4415] = 8'b00100000;
		color_arr[4416] = 8'b00100000;
		color_arr[4417] = 8'b00100000;
		color_arr[4418] = 8'b00100000;
		color_arr[4419] = 8'b00100000;
		color_arr[4420] = 8'b00100000;
		color_arr[4421] = 8'b00100000;
		color_arr[4422] = 8'b00100000;
		color_arr[4423] = 8'b00100000;
		color_arr[4424] = 8'b00100000;
		color_arr[4425] = 8'b00100000;
		color_arr[4426] = 8'b00000000;
		color_arr[4427] = 8'b00000000;
		color_arr[4428] = 8'b00000000;
		color_arr[4429] = 8'b00000000;
		color_arr[4430] = 8'b00000000;
		color_arr[4431] = 8'b00000000;
		color_arr[4432] = 8'b00000000;
		color_arr[4433] = 8'b00000000;
		color_arr[4434] = 8'b00000000;
		color_arr[4435] = 8'b00000000;
		color_arr[4436] = 8'b00000000;
		color_arr[4437] = 8'b00000000;
		color_arr[4438] = 8'b00001000;
		color_arr[4439] = 8'b00001000;
		color_arr[4440] = 8'b00001000;
		color_arr[4441] = 8'b00001000;
		color_arr[4442] = 8'b00001000;
		color_arr[4443] = 8'b00001000;
		color_arr[4444] = 8'b00001000;
		color_arr[4445] = 8'b00001000;
		color_arr[4446] = 8'b00001000;
		color_arr[4447] = 8'b00000000;
		color_arr[4448] = 8'b00000000;
		color_arr[4449] = 8'b00000000;
		color_arr[4450] = 8'b00001000;
		color_arr[4451] = 8'b00001000;
		color_arr[4452] = 8'b00001000;
		color_arr[4453] = 8'b00001000;
		color_arr[4454] = 8'b00001000;
		color_arr[4455] = 8'b00001000;
		color_arr[4456] = 8'b00001000;
		color_arr[4457] = 8'b00001000;
		color_arr[4458] = 8'b00001000;
		color_arr[4459] = 8'b00001000;
		color_arr[4460] = 8'b00001000;
		color_arr[4461] = 8'b00001000;
		color_arr[4462] = 8'b00001000;
		color_arr[4463] = 8'b00001000;
		color_arr[4464] = 8'b00001000;
		color_arr[4465] = 8'b00001000;
		color_arr[4466] = 8'b00001000;
		color_arr[4467] = 8'b00001000;
		color_arr[4468] = 8'b00001000;
		color_arr[4469] = 8'b00001000;
		color_arr[4470] = 8'b00001000;
		color_arr[4471] = 8'b00000000;
		color_arr[4472] = 8'b00000000;
		color_arr[4473] = 8'b00001000;
		color_arr[4474] = 8'b00001000;
		color_arr[4475] = 8'b00001000;
		color_arr[4476] = 8'b00001000;
		color_arr[4477] = 8'b00010010;
		color_arr[4478] = 8'b00010010;
		color_arr[4479] = 8'b00010010;
		color_arr[4480] = 8'b00010010;
		color_arr[4481] = 8'b00010010;
		color_arr[4482] = 8'b00010010;
		color_arr[4483] = 8'b00010010;
		color_arr[4484] = 8'b00010010;
		color_arr[4485] = 8'b00010010;
		color_arr[4486] = 8'b00000000;
		color_arr[4487] = 8'b00000000;
		color_arr[4488] = 8'b00000000;
		color_arr[4489] = 8'b00000010;
		color_arr[4490] = 8'b00000010;
		color_arr[4491] = 8'b00000010;
		color_arr[4492] = 8'b00000010;
		color_arr[4493] = 8'b00000010;
		color_arr[4494] = 8'b00000010;
		color_arr[4495] = 8'b00000010;
		color_arr[4496] = 8'b00000010;
		color_arr[4497] = 8'b00000010;
		color_arr[4498] = 8'b00000010;
		color_arr[4499] = 8'b00000010;
		color_arr[4500] = 8'b00000010;
		color_arr[4501] = 8'b00000010;
		color_arr[4502] = 8'b00000010;
		color_arr[4503] = 8'b00000010;
		color_arr[4504] = 8'b00000010;
		color_arr[4505] = 8'b00000010;
		color_arr[4506] = 8'b00000010;
		color_arr[4507] = 8'b00000010;
		color_arr[4508] = 8'b00000010;
		color_arr[4509] = 8'b00000010;
		color_arr[4510] = 8'b00000010;
		color_arr[4511] = 8'b00000010;
		color_arr[4512] = 8'b00000010;
		color_arr[4513] = 8'b00000010;
		color_arr[4514] = 8'b00000010;
		color_arr[4515] = 8'b00000010;
		color_arr[4516] = 8'b00000000;
		color_arr[4517] = 8'b00000000;
		color_arr[4518] = 8'b00000000;
		color_arr[4519] = 8'b00000000;
		color_arr[4520] = 8'b00000000;
		color_arr[4521] = 8'b00000000;
		color_arr[4522] = 8'b00000000;
		color_arr[4523] = 8'b00000000;
		color_arr[4524] = 8'b00100000;
		color_arr[4525] = 8'b00100000;
		color_arr[4526] = 8'b00100000;
		color_arr[4527] = 8'b00100000;
		color_arr[4528] = 8'b00100000;
		color_arr[4529] = 8'b00100000;
		color_arr[4530] = 8'b00100000;
		color_arr[4531] = 8'b00100000;
		color_arr[4532] = 8'b00100000;
		color_arr[4533] = 8'b00100000;
		color_arr[4534] = 8'b00100000;
		color_arr[4535] = 8'b00100000;
		color_arr[4536] = 8'b00100000;
		color_arr[4537] = 8'b00100000;
		color_arr[4538] = 8'b00100000;
		color_arr[4539] = 8'b00100000;
		color_arr[4540] = 8'b00100000;
		color_arr[4541] = 8'b00100000;
		color_arr[4542] = 8'b00100000;
		color_arr[4543] = 8'b00100000;
		color_arr[4544] = 8'b00100000;
		color_arr[4545] = 8'b00100000;
		color_arr[4546] = 8'b00100000;
		color_arr[4547] = 8'b00100000;
		color_arr[4548] = 8'b00100000;
		color_arr[4549] = 8'b00100000;
		color_arr[4550] = 8'b00100000;
		color_arr[4551] = 8'b00100000;
		color_arr[4552] = 8'b00100000;
		color_arr[4553] = 8'b00100000;
		color_arr[4554] = 8'b00100000;
		color_arr[4555] = 8'b00100000;
		color_arr[4556] = 8'b00100000;
		color_arr[4557] = 8'b00100000;
		color_arr[4558] = 8'b00100000;
		color_arr[4559] = 8'b00100000;
		color_arr[4560] = 8'b00000000;
		color_arr[4561] = 8'b00000000;
		color_arr[4562] = 8'b00000000;
		color_arr[4563] = 8'b00000000;
		color_arr[4564] = 8'b00000000;
		color_arr[4565] = 8'b00000000;
		color_arr[4566] = 8'b00000000;
		color_arr[4567] = 8'b00000000;
		color_arr[4568] = 8'b00000000;
		color_arr[4569] = 8'b00001000;
		color_arr[4570] = 8'b00001000;
		color_arr[4571] = 8'b00001000;
		color_arr[4572] = 8'b00001000;
		color_arr[4573] = 8'b00001000;
		color_arr[4574] = 8'b00001000;
		color_arr[4575] = 8'b00000000;
		color_arr[4576] = 8'b00000000;
		color_arr[4577] = 8'b00001000;
		color_arr[4578] = 8'b00001000;
		color_arr[4579] = 8'b00001000;
		color_arr[4580] = 8'b00001000;
		color_arr[4581] = 8'b00001000;
		color_arr[4582] = 8'b00001000;
		color_arr[4583] = 8'b00001000;
		color_arr[4584] = 8'b00001000;
		color_arr[4585] = 8'b00001000;
		color_arr[4586] = 8'b00001000;
		color_arr[4587] = 8'b00001000;
		color_arr[4588] = 8'b00001000;
		color_arr[4589] = 8'b00001000;
		color_arr[4590] = 8'b00001000;
		color_arr[4591] = 8'b00001000;
		color_arr[4592] = 8'b00001000;
		color_arr[4593] = 8'b00001000;
		color_arr[4594] = 8'b00001000;
		color_arr[4595] = 8'b00001000;
		color_arr[4596] = 8'b00001000;
		color_arr[4597] = 8'b00001000;
		color_arr[4598] = 8'b00001000;
		color_arr[4599] = 8'b00000000;
		color_arr[4600] = 8'b00000000;
		color_arr[4601] = 8'b00001000;
		color_arr[4602] = 8'b00001000;
		color_arr[4603] = 8'b00001000;
		color_arr[4604] = 8'b00001000;
		color_arr[4605] = 8'b00010010;
		color_arr[4606] = 8'b00010010;
		color_arr[4607] = 8'b00010010;
		color_arr[4608] = 8'b00010010;
		color_arr[4609] = 8'b00010010;
		color_arr[4610] = 8'b00010010;
		color_arr[4611] = 8'b00010010;
		color_arr[4612] = 8'b00010010;
		color_arr[4613] = 8'b00000000;
		color_arr[4614] = 8'b00000000;
		color_arr[4615] = 8'b00000000;
		color_arr[4616] = 8'b00000010;
		color_arr[4617] = 8'b00000010;
		color_arr[4618] = 8'b00000010;
		color_arr[4619] = 8'b00000010;
		color_arr[4620] = 8'b00000010;
		color_arr[4621] = 8'b00000010;
		color_arr[4622] = 8'b00000010;
		color_arr[4623] = 8'b00000010;
		color_arr[4624] = 8'b00000010;
		color_arr[4625] = 8'b00000010;
		color_arr[4626] = 8'b00000010;
		color_arr[4627] = 8'b00000010;
		color_arr[4628] = 8'b00000010;
		color_arr[4629] = 8'b00000010;
		color_arr[4630] = 8'b00000010;
		color_arr[4631] = 8'b00000010;
		color_arr[4632] = 8'b00000010;
		color_arr[4633] = 8'b00000010;
		color_arr[4634] = 8'b00000010;
		color_arr[4635] = 8'b00000010;
		color_arr[4636] = 8'b00000010;
		color_arr[4637] = 8'b00000010;
		color_arr[4638] = 8'b00000010;
		color_arr[4639] = 8'b00000010;
		color_arr[4640] = 8'b00000010;
		color_arr[4641] = 8'b00000010;
		color_arr[4642] = 8'b00000000;
		color_arr[4643] = 8'b00000000;
		color_arr[4644] = 8'b00000000;
		color_arr[4645] = 8'b00000000;
		color_arr[4646] = 8'b00000000;
		color_arr[4647] = 8'b00000000;
		color_arr[4648] = 8'b00100000;
		color_arr[4649] = 8'b00100000;
		color_arr[4650] = 8'b00100000;
		color_arr[4651] = 8'b00100000;
		color_arr[4652] = 8'b00100000;
		color_arr[4653] = 8'b00100000;
		color_arr[4654] = 8'b00100000;
		color_arr[4655] = 8'b00100000;
		color_arr[4656] = 8'b00100000;
		color_arr[4657] = 8'b00100000;
		color_arr[4658] = 8'b00100000;
		color_arr[4659] = 8'b00100000;
		color_arr[4660] = 8'b00100000;
		color_arr[4661] = 8'b00100000;
		color_arr[4662] = 8'b00100000;
		color_arr[4663] = 8'b00100000;
		color_arr[4664] = 8'b00100000;
		color_arr[4665] = 8'b00100000;
		color_arr[4666] = 8'b00100000;
		color_arr[4667] = 8'b00100000;
		color_arr[4668] = 8'b00100000;
		color_arr[4669] = 8'b00100000;
		color_arr[4670] = 8'b00100000;
		color_arr[4671] = 8'b00100000;
		color_arr[4672] = 8'b00100000;
		color_arr[4673] = 8'b00100000;
		color_arr[4674] = 8'b00100000;
		color_arr[4675] = 8'b00100000;
		color_arr[4676] = 8'b00100000;
		color_arr[4677] = 8'b00100000;
		color_arr[4678] = 8'b00100000;
		color_arr[4679] = 8'b00100000;
		color_arr[4680] = 8'b00100000;
		color_arr[4681] = 8'b00100000;
		color_arr[4682] = 8'b00100000;
		color_arr[4683] = 8'b00100000;
		color_arr[4684] = 8'b00100000;
		color_arr[4685] = 8'b00100000;
		color_arr[4686] = 8'b00100000;
		color_arr[4687] = 8'b00100000;
		color_arr[4688] = 8'b00001000;
		color_arr[4689] = 8'b00001000;
		color_arr[4690] = 8'b00001000;
		color_arr[4691] = 8'b00001000;
		color_arr[4692] = 8'b00001000;
		color_arr[4693] = 8'b00000000;
		color_arr[4694] = 8'b00000000;
		color_arr[4695] = 8'b00000000;
		color_arr[4696] = 8'b00000000;
		color_arr[4697] = 8'b00000000;
		color_arr[4698] = 8'b00000000;
		color_arr[4699] = 8'b00000000;
		color_arr[4700] = 8'b00001000;
		color_arr[4701] = 8'b00001000;
		color_arr[4702] = 8'b00001000;
		color_arr[4703] = 8'b00000000;
		color_arr[4704] = 8'b00000000;
		color_arr[4705] = 8'b00001000;
		color_arr[4706] = 8'b00001000;
		color_arr[4707] = 8'b00001000;
		color_arr[4708] = 8'b00001000;
		color_arr[4709] = 8'b00001000;
		color_arr[4710] = 8'b00001000;
		color_arr[4711] = 8'b00001000;
		color_arr[4712] = 8'b00001000;
		color_arr[4713] = 8'b00001000;
		color_arr[4714] = 8'b00001000;
		color_arr[4715] = 8'b00001000;
		color_arr[4716] = 8'b00001000;
		color_arr[4717] = 8'b00001000;
		color_arr[4718] = 8'b00001000;
		color_arr[4719] = 8'b00001000;
		color_arr[4720] = 8'b00001000;
		color_arr[4721] = 8'b00001000;
		color_arr[4722] = 8'b00001000;
		color_arr[4723] = 8'b00001000;
		color_arr[4724] = 8'b00001000;
		color_arr[4725] = 8'b00001000;
		color_arr[4726] = 8'b00001000;
		color_arr[4727] = 8'b00000000;
		color_arr[4728] = 8'b00000000;
		color_arr[4729] = 8'b00001000;
		color_arr[4730] = 8'b00001000;
		color_arr[4731] = 8'b00001000;
		color_arr[4732] = 8'b00001000;
		color_arr[4733] = 8'b00010010;
		color_arr[4734] = 8'b00010010;
		color_arr[4735] = 8'b00010010;
		color_arr[4736] = 8'b00010010;
		color_arr[4737] = 8'b00010010;
		color_arr[4738] = 8'b00010010;
		color_arr[4739] = 8'b00010010;
		color_arr[4740] = 8'b00010010;
		color_arr[4741] = 8'b00000000;
		color_arr[4742] = 8'b00000000;
		color_arr[4743] = 8'b00010010;
		color_arr[4744] = 8'b00000010;
		color_arr[4745] = 8'b00000010;
		color_arr[4746] = 8'b00000010;
		color_arr[4747] = 8'b00000010;
		color_arr[4748] = 8'b00000010;
		color_arr[4749] = 8'b00000010;
		color_arr[4750] = 8'b00000010;
		color_arr[4751] = 8'b00000010;
		color_arr[4752] = 8'b00000010;
		color_arr[4753] = 8'b00000010;
		color_arr[4754] = 8'b00000010;
		color_arr[4755] = 8'b00000010;
		color_arr[4756] = 8'b00000010;
		color_arr[4757] = 8'b00000010;
		color_arr[4758] = 8'b00000010;
		color_arr[4759] = 8'b00000010;
		color_arr[4760] = 8'b00000010;
		color_arr[4761] = 8'b00000010;
		color_arr[4762] = 8'b00000010;
		color_arr[4763] = 8'b00000010;
		color_arr[4764] = 8'b00000010;
		color_arr[4765] = 8'b00000010;
		color_arr[4766] = 8'b00000010;
		color_arr[4767] = 8'b00000010;
		color_arr[4768] = 8'b00000000;
		color_arr[4769] = 8'b00000000;
		color_arr[4770] = 8'b00000000;
		color_arr[4771] = 8'b00000000;
		color_arr[4772] = 8'b00000000;
		color_arr[4773] = 8'b00000010;
		color_arr[4774] = 8'b00100000;
		color_arr[4775] = 8'b00100000;
		color_arr[4776] = 8'b00100000;
		color_arr[4777] = 8'b00100000;
		color_arr[4778] = 8'b00100000;
		color_arr[4779] = 8'b00100000;
		color_arr[4780] = 8'b00100000;
		color_arr[4781] = 8'b00100000;
		color_arr[4782] = 8'b00100000;
		color_arr[4783] = 8'b00100000;
		color_arr[4784] = 8'b00100000;
		color_arr[4785] = 8'b00100000;
		color_arr[4786] = 8'b00100000;
		color_arr[4787] = 8'b00100000;
		color_arr[4788] = 8'b00100000;
		color_arr[4789] = 8'b00100000;
		color_arr[4790] = 8'b00100000;
		color_arr[4791] = 8'b00100000;
		color_arr[4792] = 8'b00100000;
		color_arr[4793] = 8'b00100000;
		color_arr[4794] = 8'b00100000;
		color_arr[4795] = 8'b00100000;
		color_arr[4796] = 8'b00100000;
		color_arr[4797] = 8'b00100000;
		color_arr[4798] = 8'b00100000;
		color_arr[4799] = 8'b00100000;
		color_arr[4800] = 8'b00100000;
		color_arr[4801] = 8'b00100000;
		color_arr[4802] = 8'b00100000;
		color_arr[4803] = 8'b00100000;
		color_arr[4804] = 8'b00100000;
		color_arr[4805] = 8'b00100000;
		color_arr[4806] = 8'b00100000;
		color_arr[4807] = 8'b00100000;
		color_arr[4808] = 8'b00100000;
		color_arr[4809] = 8'b00100000;
		color_arr[4810] = 8'b00100000;
		color_arr[4811] = 8'b00100000;
		color_arr[4812] = 8'b00100000;
		color_arr[4813] = 8'b00100000;
		color_arr[4814] = 8'b00100000;
		color_arr[4815] = 8'b00100000;
		color_arr[4816] = 8'b00001000;
		color_arr[4817] = 8'b00001000;
		color_arr[4818] = 8'b00001000;
		color_arr[4819] = 8'b00001000;
		color_arr[4820] = 8'b00001000;
		color_arr[4821] = 8'b00001000;
		color_arr[4822] = 8'b00001000;
		color_arr[4823] = 8'b00001000;
		color_arr[4824] = 8'b00000000;
		color_arr[4825] = 8'b00000000;
		color_arr[4826] = 8'b00000000;
		color_arr[4827] = 8'b00000000;
		color_arr[4828] = 8'b00000000;
		color_arr[4829] = 8'b00000000;
		color_arr[4830] = 8'b00001000;
		color_arr[4831] = 8'b00000000;
		color_arr[4832] = 8'b00000000;
		color_arr[4833] = 8'b00001000;
		color_arr[4834] = 8'b00001000;
		color_arr[4835] = 8'b00001000;
		color_arr[4836] = 8'b00001000;
		color_arr[4837] = 8'b00001000;
		color_arr[4838] = 8'b00001000;
		color_arr[4839] = 8'b00001000;
		color_arr[4840] = 8'b00001000;
		color_arr[4841] = 8'b00001000;
		color_arr[4842] = 8'b00001000;
		color_arr[4843] = 8'b00001000;
		color_arr[4844] = 8'b00001000;
		color_arr[4845] = 8'b00001000;
		color_arr[4846] = 8'b00001000;
		color_arr[4847] = 8'b00001000;
		color_arr[4848] = 8'b00001000;
		color_arr[4849] = 8'b00001000;
		color_arr[4850] = 8'b00001000;
		color_arr[4851] = 8'b00001000;
		color_arr[4852] = 8'b00001000;
		color_arr[4853] = 8'b00001000;
		color_arr[4854] = 8'b00001000;
		color_arr[4855] = 8'b00000000;
		color_arr[4856] = 8'b00000000;
		color_arr[4857] = 8'b00001000;
		color_arr[4858] = 8'b00001000;
		color_arr[4859] = 8'b00001000;
		color_arr[4860] = 8'b00001000;
		color_arr[4861] = 8'b00010010;
		color_arr[4862] = 8'b00010010;
		color_arr[4863] = 8'b00010010;
		color_arr[4864] = 8'b00010010;
		color_arr[4865] = 8'b00010010;
		color_arr[4866] = 8'b00010010;
		color_arr[4867] = 8'b00010010;
		color_arr[4868] = 8'b00000000;
		color_arr[4869] = 8'b00000000;
		color_arr[4870] = 8'b00000000;
		color_arr[4871] = 8'b00010010;
		color_arr[4872] = 8'b00000010;
		color_arr[4873] = 8'b00000010;
		color_arr[4874] = 8'b00000010;
		color_arr[4875] = 8'b00000010;
		color_arr[4876] = 8'b00000010;
		color_arr[4877] = 8'b00000010;
		color_arr[4878] = 8'b00000010;
		color_arr[4879] = 8'b00000010;
		color_arr[4880] = 8'b00000010;
		color_arr[4881] = 8'b00000010;
		color_arr[4882] = 8'b00000010;
		color_arr[4883] = 8'b00000010;
		color_arr[4884] = 8'b00000010;
		color_arr[4885] = 8'b00000010;
		color_arr[4886] = 8'b00000010;
		color_arr[4887] = 8'b00000010;
		color_arr[4888] = 8'b00000010;
		color_arr[4889] = 8'b00000010;
		color_arr[4890] = 8'b00000010;
		color_arr[4891] = 8'b00000010;
		color_arr[4892] = 8'b00000010;
		color_arr[4893] = 8'b00000010;
		color_arr[4894] = 8'b00000010;
		color_arr[4895] = 8'b00000000;
		color_arr[4896] = 8'b00000000;
		color_arr[4897] = 8'b00000000;
		color_arr[4898] = 8'b00000000;
		color_arr[4899] = 8'b00000010;
		color_arr[4900] = 8'b00000010;
		color_arr[4901] = 8'b00000010;
		color_arr[4902] = 8'b00100000;
		color_arr[4903] = 8'b00100000;
		color_arr[4904] = 8'b00100000;
		color_arr[4905] = 8'b00100000;
		color_arr[4906] = 8'b00100000;
		color_arr[4907] = 8'b00100000;
		color_arr[4908] = 8'b00100000;
		color_arr[4909] = 8'b00100000;
		color_arr[4910] = 8'b00100000;
		color_arr[4911] = 8'b00100000;
		color_arr[4912] = 8'b00100000;
		color_arr[4913] = 8'b00100000;
		color_arr[4914] = 8'b00100000;
		color_arr[4915] = 8'b00100000;
		color_arr[4916] = 8'b00100000;
		color_arr[4917] = 8'b00100000;
		color_arr[4918] = 8'b00100000;
		color_arr[4919] = 8'b00100000;
		color_arr[4920] = 8'b00100000;
		color_arr[4921] = 8'b00100000;
		color_arr[4922] = 8'b00100000;
		color_arr[4923] = 8'b00100000;
		color_arr[4924] = 8'b00100000;
		color_arr[4925] = 8'b00100000;
		color_arr[4926] = 8'b00100000;
		color_arr[4927] = 8'b00100000;
		color_arr[4928] = 8'b00100000;
		color_arr[4929] = 8'b00100000;
		color_arr[4930] = 8'b00100000;
		color_arr[4931] = 8'b00100000;
		color_arr[4932] = 8'b00100000;
		color_arr[4933] = 8'b00100000;
		color_arr[4934] = 8'b00100000;
		color_arr[4935] = 8'b00100000;
		color_arr[4936] = 8'b00100000;
		color_arr[4937] = 8'b00100000;
		color_arr[4938] = 8'b00100000;
		color_arr[4939] = 8'b00100000;
		color_arr[4940] = 8'b00100000;
		color_arr[4941] = 8'b00100000;
		color_arr[4942] = 8'b00100000;
		color_arr[4943] = 8'b00100000;
		color_arr[4944] = 8'b00001000;
		color_arr[4945] = 8'b00001000;
		color_arr[4946] = 8'b00001000;
		color_arr[4947] = 8'b00001000;
		color_arr[4948] = 8'b00001000;
		color_arr[4949] = 8'b00001000;
		color_arr[4950] = 8'b00001000;
		color_arr[4951] = 8'b00001000;
		color_arr[4952] = 8'b00001000;
		color_arr[4953] = 8'b00001000;
		color_arr[4954] = 8'b00001000;
		color_arr[4955] = 8'b00000000;
		color_arr[4956] = 8'b00000000;
		color_arr[4957] = 8'b00000000;
		color_arr[4958] = 8'b00000000;
		color_arr[4959] = 8'b00000000;
		color_arr[4960] = 8'b00000000;
		color_arr[4961] = 8'b00001000;
		color_arr[4962] = 8'b00001000;
		color_arr[4963] = 8'b00001000;
		color_arr[4964] = 8'b00001000;
		color_arr[4965] = 8'b00001000;
		color_arr[4966] = 8'b00001000;
		color_arr[4967] = 8'b00001000;
		color_arr[4968] = 8'b00001000;
		color_arr[4969] = 8'b00001000;
		color_arr[4970] = 8'b00001000;
		color_arr[4971] = 8'b00001000;
		color_arr[4972] = 8'b00001000;
		color_arr[4973] = 8'b00001000;
		color_arr[4974] = 8'b00001000;
		color_arr[4975] = 8'b00001000;
		color_arr[4976] = 8'b00001000;
		color_arr[4977] = 8'b00001000;
		color_arr[4978] = 8'b00001000;
		color_arr[4979] = 8'b00001000;
		color_arr[4980] = 8'b00001000;
		color_arr[4981] = 8'b00001000;
		color_arr[4982] = 8'b00001000;
		color_arr[4983] = 8'b00000000;
		color_arr[4984] = 8'b00000000;
		color_arr[4985] = 8'b00001000;
		color_arr[4986] = 8'b00001000;
		color_arr[4987] = 8'b00001000;
		color_arr[4988] = 8'b00001000;
		color_arr[4989] = 8'b00010010;
		color_arr[4990] = 8'b00010010;
		color_arr[4991] = 8'b00010010;
		color_arr[4992] = 8'b00010010;
		color_arr[4993] = 8'b00010010;
		color_arr[4994] = 8'b00010010;
		color_arr[4995] = 8'b00010010;
		color_arr[4996] = 8'b00000000;
		color_arr[4997] = 8'b00000000;
		color_arr[4998] = 8'b00010010;
		color_arr[4999] = 8'b00010010;
		color_arr[5000] = 8'b00000010;
		color_arr[5001] = 8'b00000010;
		color_arr[5002] = 8'b00000010;
		color_arr[5003] = 8'b00000010;
		color_arr[5004] = 8'b00000010;
		color_arr[5005] = 8'b00000010;
		color_arr[5006] = 8'b00000010;
		color_arr[5007] = 8'b00000010;
		color_arr[5008] = 8'b00000010;
		color_arr[5009] = 8'b00000010;
		color_arr[5010] = 8'b00000010;
		color_arr[5011] = 8'b00000010;
		color_arr[5012] = 8'b00000010;
		color_arr[5013] = 8'b00000010;
		color_arr[5014] = 8'b00000010;
		color_arr[5015] = 8'b00000010;
		color_arr[5016] = 8'b00000010;
		color_arr[5017] = 8'b00000010;
		color_arr[5018] = 8'b00000010;
		color_arr[5019] = 8'b00000010;
		color_arr[5020] = 8'b00000010;
		color_arr[5021] = 8'b00000010;
		color_arr[5022] = 8'b00000000;
		color_arr[5023] = 8'b00000000;
		color_arr[5024] = 8'b00000000;
		color_arr[5025] = 8'b00000010;
		color_arr[5026] = 8'b00000010;
		color_arr[5027] = 8'b00000010;
		color_arr[5028] = 8'b00000010;
		color_arr[5029] = 8'b00000010;
		color_arr[5030] = 8'b00100000;
		color_arr[5031] = 8'b00100000;
		color_arr[5032] = 8'b00100000;
		color_arr[5033] = 8'b00100000;
		color_arr[5034] = 8'b00100000;
		color_arr[5035] = 8'b00100000;
		color_arr[5036] = 8'b00100000;
		color_arr[5037] = 8'b00100000;
		color_arr[5038] = 8'b00100000;
		color_arr[5039] = 8'b00100000;
		color_arr[5040] = 8'b00100000;
		color_arr[5041] = 8'b00100000;
		color_arr[5042] = 8'b00100000;
		color_arr[5043] = 8'b00100000;
		color_arr[5044] = 8'b00100000;
		color_arr[5045] = 8'b00100000;
		color_arr[5046] = 8'b00100000;
		color_arr[5047] = 8'b00100000;
		color_arr[5048] = 8'b00100000;
		color_arr[5049] = 8'b00100000;
		color_arr[5050] = 8'b00100000;
		color_arr[5051] = 8'b00100000;
		color_arr[5052] = 8'b00100000;
		color_arr[5053] = 8'b00100000;
		color_arr[5054] = 8'b00100000;
		color_arr[5055] = 8'b00100000;
		color_arr[5056] = 8'b00100000;
		color_arr[5057] = 8'b00100000;
		color_arr[5058] = 8'b00100000;
		color_arr[5059] = 8'b00100000;
		color_arr[5060] = 8'b00100000;
		color_arr[5061] = 8'b00100000;
		color_arr[5062] = 8'b00100000;
		color_arr[5063] = 8'b00100000;
		color_arr[5064] = 8'b00100000;
		color_arr[5065] = 8'b00100000;
		color_arr[5066] = 8'b00100000;
		color_arr[5067] = 8'b00100000;
		color_arr[5068] = 8'b00100000;
		color_arr[5069] = 8'b00100000;
		color_arr[5070] = 8'b00100000;
		color_arr[5071] = 8'b00100000;
		color_arr[5072] = 8'b00001000;
		color_arr[5073] = 8'b00001000;
		color_arr[5074] = 8'b00001000;
		color_arr[5075] = 8'b00001000;
		color_arr[5076] = 8'b00001000;
		color_arr[5077] = 8'b00001000;
		color_arr[5078] = 8'b00001000;
		color_arr[5079] = 8'b00001000;
		color_arr[5080] = 8'b00001000;
		color_arr[5081] = 8'b00001000;
		color_arr[5082] = 8'b00001000;
		color_arr[5083] = 8'b00001000;
		color_arr[5084] = 8'b00001000;
		color_arr[5085] = 8'b00000000;
		color_arr[5086] = 8'b00000000;
		color_arr[5087] = 8'b00000000;
		color_arr[5088] = 8'b00000000;
		color_arr[5089] = 8'b00001000;
		color_arr[5090] = 8'b00001000;
		color_arr[5091] = 8'b00001000;
		color_arr[5092] = 8'b00001000;
		color_arr[5093] = 8'b00001000;
		color_arr[5094] = 8'b00001000;
		color_arr[5095] = 8'b00001000;
		color_arr[5096] = 8'b00001000;
		color_arr[5097] = 8'b00001000;
		color_arr[5098] = 8'b00001000;
		color_arr[5099] = 8'b00001000;
		color_arr[5100] = 8'b00001000;
		color_arr[5101] = 8'b00001000;
		color_arr[5102] = 8'b00001000;
		color_arr[5103] = 8'b00001000;
		color_arr[5104] = 8'b00001000;
		color_arr[5105] = 8'b00001000;
		color_arr[5106] = 8'b00001000;
		color_arr[5107] = 8'b00001000;
		color_arr[5108] = 8'b00001000;
		color_arr[5109] = 8'b00001000;
		color_arr[5110] = 8'b00000000;
		color_arr[5111] = 8'b00000000;
		color_arr[5112] = 8'b00000000;
		color_arr[5113] = 8'b00001000;
		color_arr[5114] = 8'b00001000;
		color_arr[5115] = 8'b00001000;
		color_arr[5116] = 8'b00001000;
		color_arr[5117] = 8'b00010010;
		color_arr[5118] = 8'b00010010;
		color_arr[5119] = 8'b00010010;
		color_arr[5120] = 8'b00010010;
		color_arr[5121] = 8'b00010010;
		color_arr[5122] = 8'b00010010;
		color_arr[5123] = 8'b00000000;
		color_arr[5124] = 8'b00000000;
		color_arr[5125] = 8'b00000000;
		color_arr[5126] = 8'b00010010;
		color_arr[5127] = 8'b00010010;
		color_arr[5128] = 8'b00000010;
		color_arr[5129] = 8'b00000010;
		color_arr[5130] = 8'b00000010;
		color_arr[5131] = 8'b00000010;
		color_arr[5132] = 8'b00000010;
		color_arr[5133] = 8'b00000010;
		color_arr[5134] = 8'b00000010;
		color_arr[5135] = 8'b00000010;
		color_arr[5136] = 8'b00000010;
		color_arr[5137] = 8'b00000010;
		color_arr[5138] = 8'b00000010;
		color_arr[5139] = 8'b00000010;
		color_arr[5140] = 8'b00000010;
		color_arr[5141] = 8'b00000010;
		color_arr[5142] = 8'b00000010;
		color_arr[5143] = 8'b00000010;
		color_arr[5144] = 8'b00000010;
		color_arr[5145] = 8'b00000010;
		color_arr[5146] = 8'b00000010;
		color_arr[5147] = 8'b00000010;
		color_arr[5148] = 8'b00000000;
		color_arr[5149] = 8'b00000000;
		color_arr[5150] = 8'b00000000;
		color_arr[5151] = 8'b00000000;
		color_arr[5152] = 8'b00000010;
		color_arr[5153] = 8'b00000010;
		color_arr[5154] = 8'b00000010;
		color_arr[5155] = 8'b00000010;
		color_arr[5156] = 8'b00000010;
		color_arr[5157] = 8'b00000010;
		color_arr[5158] = 8'b00100000;
		color_arr[5159] = 8'b00100000;
		color_arr[5160] = 8'b00100000;
		color_arr[5161] = 8'b00100000;
		color_arr[5162] = 8'b00100000;
		color_arr[5163] = 8'b00100000;
		color_arr[5164] = 8'b00100000;
		color_arr[5165] = 8'b00100000;
		color_arr[5166] = 8'b00100000;
		color_arr[5167] = 8'b00100000;
		color_arr[5168] = 8'b00100000;
		color_arr[5169] = 8'b00100000;
		color_arr[5170] = 8'b00100000;
		color_arr[5171] = 8'b00100000;
		color_arr[5172] = 8'b00100000;
		color_arr[5173] = 8'b00100000;
		color_arr[5174] = 8'b00100000;
		color_arr[5175] = 8'b00100000;
		color_arr[5176] = 8'b00100000;
		color_arr[5177] = 8'b00100000;
		color_arr[5178] = 8'b00100000;
		color_arr[5179] = 8'b00100000;
		color_arr[5180] = 8'b00100000;
		color_arr[5181] = 8'b00100000;
		color_arr[5182] = 8'b00100000;
		color_arr[5183] = 8'b00100000;
		color_arr[5184] = 8'b00100000;
		color_arr[5185] = 8'b00100000;
		color_arr[5186] = 8'b00100000;
		color_arr[5187] = 8'b00100000;
		color_arr[5188] = 8'b00100000;
		color_arr[5189] = 8'b00100000;
		color_arr[5190] = 8'b00100000;
		color_arr[5191] = 8'b00100000;
		color_arr[5192] = 8'b00100000;
		color_arr[5193] = 8'b00100000;
		color_arr[5194] = 8'b00100000;
		color_arr[5195] = 8'b00100000;
		color_arr[5196] = 8'b00100000;
		color_arr[5197] = 8'b00100000;
		color_arr[5198] = 8'b00100000;
		color_arr[5199] = 8'b00100000;
		color_arr[5200] = 8'b00001000;
		color_arr[5201] = 8'b00001000;
		color_arr[5202] = 8'b00001000;
		color_arr[5203] = 8'b00001000;
		color_arr[5204] = 8'b00001000;
		color_arr[5205] = 8'b00001000;
		color_arr[5206] = 8'b00001000;
		color_arr[5207] = 8'b00001000;
		color_arr[5208] = 8'b00001000;
		color_arr[5209] = 8'b00001000;
		color_arr[5210] = 8'b00001000;
		color_arr[5211] = 8'b00001000;
		color_arr[5212] = 8'b00001000;
		color_arr[5213] = 8'b00001000;
		color_arr[5214] = 8'b00000000;
		color_arr[5215] = 8'b00000000;
		color_arr[5216] = 8'b00000000;
		color_arr[5217] = 8'b00000000;
		color_arr[5218] = 8'b00001000;
		color_arr[5219] = 8'b00001000;
		color_arr[5220] = 8'b00001000;
		color_arr[5221] = 8'b00001000;
		color_arr[5222] = 8'b00001000;
		color_arr[5223] = 8'b00001000;
		color_arr[5224] = 8'b00001000;
		color_arr[5225] = 8'b00001000;
		color_arr[5226] = 8'b00001000;
		color_arr[5227] = 8'b00001000;
		color_arr[5228] = 8'b00001000;
		color_arr[5229] = 8'b00001000;
		color_arr[5230] = 8'b00001000;
		color_arr[5231] = 8'b00001000;
		color_arr[5232] = 8'b00001000;
		color_arr[5233] = 8'b00001000;
		color_arr[5234] = 8'b00001000;
		color_arr[5235] = 8'b00001000;
		color_arr[5236] = 8'b00001000;
		color_arr[5237] = 8'b00001000;
		color_arr[5238] = 8'b00000000;
		color_arr[5239] = 8'b00000000;
		color_arr[5240] = 8'b00001000;
		color_arr[5241] = 8'b00001000;
		color_arr[5242] = 8'b00001000;
		color_arr[5243] = 8'b00001000;
		color_arr[5244] = 8'b00001000;
		color_arr[5245] = 8'b00010010;
		color_arr[5246] = 8'b00010010;
		color_arr[5247] = 8'b00010010;
		color_arr[5248] = 8'b00010010;
		color_arr[5249] = 8'b00010010;
		color_arr[5250] = 8'b00010010;
		color_arr[5251] = 8'b00000000;
		color_arr[5252] = 8'b00000000;
		color_arr[5253] = 8'b00010010;
		color_arr[5254] = 8'b00010010;
		color_arr[5255] = 8'b00010010;
		color_arr[5256] = 8'b00000010;
		color_arr[5257] = 8'b00000010;
		color_arr[5258] = 8'b00000010;
		color_arr[5259] = 8'b00000010;
		color_arr[5260] = 8'b00000010;
		color_arr[5261] = 8'b00000010;
		color_arr[5262] = 8'b00000010;
		color_arr[5263] = 8'b00000010;
		color_arr[5264] = 8'b00000010;
		color_arr[5265] = 8'b00000010;
		color_arr[5266] = 8'b00000010;
		color_arr[5267] = 8'b00000010;
		color_arr[5268] = 8'b00000010;
		color_arr[5269] = 8'b00000010;
		color_arr[5270] = 8'b00000010;
		color_arr[5271] = 8'b00000010;
		color_arr[5272] = 8'b00000010;
		color_arr[5273] = 8'b00000010;
		color_arr[5274] = 8'b00000010;
		color_arr[5275] = 8'b00000000;
		color_arr[5276] = 8'b00000000;
		color_arr[5277] = 8'b00000000;
		color_arr[5278] = 8'b00000000;
		color_arr[5279] = 8'b00000010;
		color_arr[5280] = 8'b00000010;
		color_arr[5281] = 8'b00000010;
		color_arr[5282] = 8'b00000010;
		color_arr[5283] = 8'b00000010;
		color_arr[5284] = 8'b00000010;
		color_arr[5285] = 8'b00000010;
		color_arr[5286] = 8'b00100000;
		color_arr[5287] = 8'b00100000;
		color_arr[5288] = 8'b00100000;
		color_arr[5289] = 8'b00100000;
		color_arr[5290] = 8'b00100000;
		color_arr[5291] = 8'b00100000;
		color_arr[5292] = 8'b00100000;
		color_arr[5293] = 8'b00100000;
		color_arr[5294] = 8'b00100000;
		color_arr[5295] = 8'b00100000;
		color_arr[5296] = 8'b00100000;
		color_arr[5297] = 8'b00100000;
		color_arr[5298] = 8'b00100000;
		color_arr[5299] = 8'b00100000;
		color_arr[5300] = 8'b00100000;
		color_arr[5301] = 8'b00100000;
		color_arr[5302] = 8'b00100000;
		color_arr[5303] = 8'b00100000;
		color_arr[5304] = 8'b00100000;
		color_arr[5305] = 8'b00100000;
		color_arr[5306] = 8'b00100000;
		color_arr[5307] = 8'b00100000;
		color_arr[5308] = 8'b00100000;
		color_arr[5309] = 8'b00100000;
		color_arr[5310] = 8'b00100000;
		color_arr[5311] = 8'b00100000;
		color_arr[5312] = 8'b00100000;
		color_arr[5313] = 8'b00100000;
		color_arr[5314] = 8'b00100000;
		color_arr[5315] = 8'b00100000;
		color_arr[5316] = 8'b00100000;
		color_arr[5317] = 8'b00100000;
		color_arr[5318] = 8'b00100000;
		color_arr[5319] = 8'b00100000;
		color_arr[5320] = 8'b00100000;
		color_arr[5321] = 8'b00100000;
		color_arr[5322] = 8'b00100000;
		color_arr[5323] = 8'b00100000;
		color_arr[5324] = 8'b00100000;
		color_arr[5325] = 8'b00100000;
		color_arr[5326] = 8'b00100000;
		color_arr[5327] = 8'b00100000;
		color_arr[5328] = 8'b00001000;
		color_arr[5329] = 8'b00001000;
		color_arr[5330] = 8'b00001000;
		color_arr[5331] = 8'b00001000;
		color_arr[5332] = 8'b00001000;
		color_arr[5333] = 8'b00001000;
		color_arr[5334] = 8'b00001000;
		color_arr[5335] = 8'b00001000;
		color_arr[5336] = 8'b00001000;
		color_arr[5337] = 8'b00001000;
		color_arr[5338] = 8'b00001000;
		color_arr[5339] = 8'b00001000;
		color_arr[5340] = 8'b00001000;
		color_arr[5341] = 8'b00001000;
		color_arr[5342] = 8'b00001000;
		color_arr[5343] = 8'b00001000;
		color_arr[5344] = 8'b00000000;
		color_arr[5345] = 8'b00000000;
		color_arr[5346] = 8'b00000000;
		color_arr[5347] = 8'b00001000;
		color_arr[5348] = 8'b00001000;
		color_arr[5349] = 8'b00001000;
		color_arr[5350] = 8'b00001000;
		color_arr[5351] = 8'b00001000;
		color_arr[5352] = 8'b00001000;
		color_arr[5353] = 8'b00001000;
		color_arr[5354] = 8'b00001000;
		color_arr[5355] = 8'b00001000;
		color_arr[5356] = 8'b00001000;
		color_arr[5357] = 8'b00001000;
		color_arr[5358] = 8'b00001000;
		color_arr[5359] = 8'b00001000;
		color_arr[5360] = 8'b00001000;
		color_arr[5361] = 8'b00001000;
		color_arr[5362] = 8'b00001000;
		color_arr[5363] = 8'b00001000;
		color_arr[5364] = 8'b00001000;
		color_arr[5365] = 8'b00000000;
		color_arr[5366] = 8'b00000000;
		color_arr[5367] = 8'b00000000;
		color_arr[5368] = 8'b00001000;
		color_arr[5369] = 8'b00001000;
		color_arr[5370] = 8'b00001000;
		color_arr[5371] = 8'b00001000;
		color_arr[5372] = 8'b00001000;
		color_arr[5373] = 8'b00010010;
		color_arr[5374] = 8'b00010010;
		color_arr[5375] = 8'b00010010;
		color_arr[5376] = 8'b00010010;
		color_arr[5377] = 8'b00010010;
		color_arr[5378] = 8'b00010010;
		color_arr[5379] = 8'b00000000;
		color_arr[5380] = 8'b00000000;
		color_arr[5381] = 8'b00010010;
		color_arr[5382] = 8'b00010010;
		color_arr[5383] = 8'b00010010;
		color_arr[5384] = 8'b00000010;
		color_arr[5385] = 8'b00000010;
		color_arr[5386] = 8'b00000010;
		color_arr[5387] = 8'b00000010;
		color_arr[5388] = 8'b00000010;
		color_arr[5389] = 8'b00000010;
		color_arr[5390] = 8'b00000010;
		color_arr[5391] = 8'b00000010;
		color_arr[5392] = 8'b00000010;
		color_arr[5393] = 8'b00000010;
		color_arr[5394] = 8'b00000010;
		color_arr[5395] = 8'b00000010;
		color_arr[5396] = 8'b00000010;
		color_arr[5397] = 8'b00000010;
		color_arr[5398] = 8'b00000010;
		color_arr[5399] = 8'b00000010;
		color_arr[5400] = 8'b00000010;
		color_arr[5401] = 8'b00000010;
		color_arr[5402] = 8'b00000000;
		color_arr[5403] = 8'b00000000;
		color_arr[5404] = 8'b00000000;
		color_arr[5405] = 8'b00000010;
		color_arr[5406] = 8'b00000010;
		color_arr[5407] = 8'b00000010;
		color_arr[5408] = 8'b00000010;
		color_arr[5409] = 8'b00000010;
		color_arr[5410] = 8'b00000010;
		color_arr[5411] = 8'b00000010;
		color_arr[5412] = 8'b00000010;
		color_arr[5413] = 8'b00000010;
		color_arr[5414] = 8'b00100000;
		color_arr[5415] = 8'b00100000;
		color_arr[5416] = 8'b00100000;
		color_arr[5417] = 8'b00100000;
		color_arr[5418] = 8'b00100000;
		color_arr[5419] = 8'b00100000;
		color_arr[5420] = 8'b00100000;
		color_arr[5421] = 8'b00100000;
		color_arr[5422] = 8'b00100000;
		color_arr[5423] = 8'b00100000;
		color_arr[5424] = 8'b00100000;
		color_arr[5425] = 8'b00100000;
		color_arr[5426] = 8'b00100000;
		color_arr[5427] = 8'b00100000;
		color_arr[5428] = 8'b00100000;
		color_arr[5429] = 8'b00100000;
		color_arr[5430] = 8'b00100000;
		color_arr[5431] = 8'b00100000;
		color_arr[5432] = 8'b00100000;
		color_arr[5433] = 8'b00100000;
		color_arr[5434] = 8'b00100000;
		color_arr[5435] = 8'b00100000;
		color_arr[5436] = 8'b00100000;
		color_arr[5437] = 8'b00100000;
		color_arr[5438] = 8'b00100000;
		color_arr[5439] = 8'b00100000;
		color_arr[5440] = 8'b00100000;
		color_arr[5441] = 8'b00100000;
		color_arr[5442] = 8'b00100000;
		color_arr[5443] = 8'b00100000;
		color_arr[5444] = 8'b00100000;
		color_arr[5445] = 8'b00100000;
		color_arr[5446] = 8'b00100000;
		color_arr[5447] = 8'b00100000;
		color_arr[5448] = 8'b00100000;
		color_arr[5449] = 8'b00100000;
		color_arr[5450] = 8'b00100000;
		color_arr[5451] = 8'b00100000;
		color_arr[5452] = 8'b00100000;
		color_arr[5453] = 8'b00100000;
		color_arr[5454] = 8'b00100000;
		color_arr[5455] = 8'b00100000;
		color_arr[5456] = 8'b00001000;
		color_arr[5457] = 8'b00001000;
		color_arr[5458] = 8'b00001000;
		color_arr[5459] = 8'b00001000;
		color_arr[5460] = 8'b00001000;
		color_arr[5461] = 8'b00001000;
		color_arr[5462] = 8'b00001000;
		color_arr[5463] = 8'b00001000;
		color_arr[5464] = 8'b00001000;
		color_arr[5465] = 8'b00001000;
		color_arr[5466] = 8'b00001000;
		color_arr[5467] = 8'b00001000;
		color_arr[5468] = 8'b00001000;
		color_arr[5469] = 8'b00001000;
		color_arr[5470] = 8'b00001000;
		color_arr[5471] = 8'b00001000;
		color_arr[5472] = 8'b00000000;
		color_arr[5473] = 8'b00000000;
		color_arr[5474] = 8'b00000000;
		color_arr[5475] = 8'b00001000;
		color_arr[5476] = 8'b00001000;
		color_arr[5477] = 8'b00001000;
		color_arr[5478] = 8'b00001000;
		color_arr[5479] = 8'b00001000;
		color_arr[5480] = 8'b00001000;
		color_arr[5481] = 8'b00001000;
		color_arr[5482] = 8'b00001000;
		color_arr[5483] = 8'b00001000;
		color_arr[5484] = 8'b00001000;
		color_arr[5485] = 8'b00001000;
		color_arr[5486] = 8'b00001000;
		color_arr[5487] = 8'b00001000;
		color_arr[5488] = 8'b00001000;
		color_arr[5489] = 8'b00001000;
		color_arr[5490] = 8'b00001000;
		color_arr[5491] = 8'b00001000;
		color_arr[5492] = 8'b00001000;
		color_arr[5493] = 8'b00000000;
		color_arr[5494] = 8'b00000000;
		color_arr[5495] = 8'b00001000;
		color_arr[5496] = 8'b00001000;
		color_arr[5497] = 8'b00001000;
		color_arr[5498] = 8'b00001000;
		color_arr[5499] = 8'b00001000;
		color_arr[5500] = 8'b00001000;
		color_arr[5501] = 8'b00010010;
		color_arr[5502] = 8'b00010010;
		color_arr[5503] = 8'b00010010;
		color_arr[5504] = 8'b00010010;
		color_arr[5505] = 8'b00010010;
		color_arr[5506] = 8'b00010010;
		color_arr[5507] = 8'b00000000;
		color_arr[5508] = 8'b00000000;
		color_arr[5509] = 8'b00010010;
		color_arr[5510] = 8'b00010010;
		color_arr[5511] = 8'b00010010;
		color_arr[5512] = 8'b00000010;
		color_arr[5513] = 8'b00000010;
		color_arr[5514] = 8'b00000010;
		color_arr[5515] = 8'b00000010;
		color_arr[5516] = 8'b00000010;
		color_arr[5517] = 8'b00000010;
		color_arr[5518] = 8'b00000010;
		color_arr[5519] = 8'b00000010;
		color_arr[5520] = 8'b00000010;
		color_arr[5521] = 8'b00000010;
		color_arr[5522] = 8'b00000010;
		color_arr[5523] = 8'b00000010;
		color_arr[5524] = 8'b00000010;
		color_arr[5525] = 8'b00000010;
		color_arr[5526] = 8'b00000010;
		color_arr[5527] = 8'b00000010;
		color_arr[5528] = 8'b00000010;
		color_arr[5529] = 8'b00000010;
		color_arr[5530] = 8'b00000000;
		color_arr[5531] = 8'b00000000;
		color_arr[5532] = 8'b00000010;
		color_arr[5533] = 8'b00000010;
		color_arr[5534] = 8'b00000010;
		color_arr[5535] = 8'b00000010;
		color_arr[5536] = 8'b00000010;
		color_arr[5537] = 8'b00000010;
		color_arr[5538] = 8'b00000010;
		color_arr[5539] = 8'b00000010;
		color_arr[5540] = 8'b00000010;
		color_arr[5541] = 8'b00000010;
		color_arr[5542] = 8'b00100000;
		color_arr[5543] = 8'b00100000;
		color_arr[5544] = 8'b00100000;
		color_arr[5545] = 8'b00100000;
		color_arr[5546] = 8'b00100000;
		color_arr[5547] = 8'b00100000;
		color_arr[5548] = 8'b00100000;
		color_arr[5549] = 8'b00100000;
		color_arr[5550] = 8'b00100000;
		color_arr[5551] = 8'b00100000;
		color_arr[5552] = 8'b00100000;
		color_arr[5553] = 8'b00100000;
		color_arr[5554] = 8'b00100000;
		color_arr[5555] = 8'b00100000;
		color_arr[5556] = 8'b00100000;
		color_arr[5557] = 8'b00100000;
		color_arr[5558] = 8'b00100000;
		color_arr[5559] = 8'b00100000;
		color_arr[5560] = 8'b00100000;
		color_arr[5561] = 8'b00100000;
		color_arr[5562] = 8'b00100000;
		color_arr[5563] = 8'b00100000;
		color_arr[5564] = 8'b00100000;
		color_arr[5565] = 8'b00100000;
		color_arr[5566] = 8'b00100000;
		color_arr[5567] = 8'b00100000;
		color_arr[5568] = 8'b00100000;
		color_arr[5569] = 8'b00100000;
		color_arr[5570] = 8'b00100000;
		color_arr[5571] = 8'b00100000;
		color_arr[5572] = 8'b00100000;
		color_arr[5573] = 8'b00100000;
		color_arr[5574] = 8'b00100000;
		color_arr[5575] = 8'b00100000;
		color_arr[5576] = 8'b00100000;
		color_arr[5577] = 8'b00100000;
		color_arr[5578] = 8'b00100000;
		color_arr[5579] = 8'b00100000;
		color_arr[5580] = 8'b00100000;
		color_arr[5581] = 8'b00100000;
		color_arr[5582] = 8'b00100000;
		color_arr[5583] = 8'b00100000;
		color_arr[5584] = 8'b00001000;
		color_arr[5585] = 8'b00001000;
		color_arr[5586] = 8'b00001000;
		color_arr[5587] = 8'b00001000;
		color_arr[5588] = 8'b00001000;
		color_arr[5589] = 8'b00001000;
		color_arr[5590] = 8'b00001000;
		color_arr[5591] = 8'b00001000;
		color_arr[5592] = 8'b00001000;
		color_arr[5593] = 8'b00001000;
		color_arr[5594] = 8'b00001000;
		color_arr[5595] = 8'b00001000;
		color_arr[5596] = 8'b00001000;
		color_arr[5597] = 8'b00001000;
		color_arr[5598] = 8'b00001000;
		color_arr[5599] = 8'b00001000;
		color_arr[5600] = 8'b00001000;
		color_arr[5601] = 8'b00000000;
		color_arr[5602] = 8'b00000000;
		color_arr[5603] = 8'b00000000;
		color_arr[5604] = 8'b00001000;
		color_arr[5605] = 8'b00001000;
		color_arr[5606] = 8'b00001000;
		color_arr[5607] = 8'b00001000;
		color_arr[5608] = 8'b00001000;
		color_arr[5609] = 8'b00001000;
		color_arr[5610] = 8'b00001000;
		color_arr[5611] = 8'b00001000;
		color_arr[5612] = 8'b00001000;
		color_arr[5613] = 8'b00001000;
		color_arr[5614] = 8'b00001000;
		color_arr[5615] = 8'b00001000;
		color_arr[5616] = 8'b00001000;
		color_arr[5617] = 8'b00001000;
		color_arr[5618] = 8'b00001000;
		color_arr[5619] = 8'b00001000;
		color_arr[5620] = 8'b00001000;
		color_arr[5621] = 8'b00000000;
		color_arr[5622] = 8'b00000000;
		color_arr[5623] = 8'b00001000;
		color_arr[5624] = 8'b00001000;
		color_arr[5625] = 8'b00001000;
		color_arr[5626] = 8'b00001000;
		color_arr[5627] = 8'b00001000;
		color_arr[5628] = 8'b00001000;
		color_arr[5629] = 8'b00010010;
		color_arr[5630] = 8'b00010010;
		color_arr[5631] = 8'b00010010;
		color_arr[5632] = 8'b00010010;
		color_arr[5633] = 8'b00010010;
		color_arr[5634] = 8'b00000000;
		color_arr[5635] = 8'b00000000;
		color_arr[5636] = 8'b00000000;
		color_arr[5637] = 8'b00010010;
		color_arr[5638] = 8'b00010010;
		color_arr[5639] = 8'b00010010;
		color_arr[5640] = 8'b00000010;
		color_arr[5641] = 8'b00000010;
		color_arr[5642] = 8'b00000010;
		color_arr[5643] = 8'b00000010;
		color_arr[5644] = 8'b00000010;
		color_arr[5645] = 8'b00000010;
		color_arr[5646] = 8'b00000010;
		color_arr[5647] = 8'b00000010;
		color_arr[5648] = 8'b00000010;
		color_arr[5649] = 8'b00000010;
		color_arr[5650] = 8'b00000010;
		color_arr[5651] = 8'b00000010;
		color_arr[5652] = 8'b00000010;
		color_arr[5653] = 8'b00000010;
		color_arr[5654] = 8'b00000010;
		color_arr[5655] = 8'b00000010;
		color_arr[5656] = 8'b00000010;
		color_arr[5657] = 8'b00000000;
		color_arr[5658] = 8'b00000000;
		color_arr[5659] = 8'b00000000;
		color_arr[5660] = 8'b00000010;
		color_arr[5661] = 8'b00000010;
		color_arr[5662] = 8'b00000010;
		color_arr[5663] = 8'b00000010;
		color_arr[5664] = 8'b00000010;
		color_arr[5665] = 8'b00000010;
		color_arr[5666] = 8'b00000010;
		color_arr[5667] = 8'b00000010;
		color_arr[5668] = 8'b00000010;
		color_arr[5669] = 8'b00000010;
		color_arr[5670] = 8'b00100000;
		color_arr[5671] = 8'b00100000;
		color_arr[5672] = 8'b00100000;
		color_arr[5673] = 8'b00100000;
		color_arr[5674] = 8'b00100000;
		color_arr[5675] = 8'b00100000;
		color_arr[5676] = 8'b00100000;
		color_arr[5677] = 8'b00100000;
		color_arr[5678] = 8'b00100000;
		color_arr[5679] = 8'b00100000;
		color_arr[5680] = 8'b00100000;
		color_arr[5681] = 8'b00100000;
		color_arr[5682] = 8'b00100000;
		color_arr[5683] = 8'b00100000;
		color_arr[5684] = 8'b00100000;
		color_arr[5685] = 8'b00100000;
		color_arr[5686] = 8'b00100000;
		color_arr[5687] = 8'b00100000;
		color_arr[5688] = 8'b00100000;
		color_arr[5689] = 8'b00100000;
		color_arr[5690] = 8'b00100000;
		color_arr[5691] = 8'b00100000;
		color_arr[5692] = 8'b00100000;
		color_arr[5693] = 8'b00100000;
		color_arr[5694] = 8'b00100000;
		color_arr[5695] = 8'b00100000;
		color_arr[5696] = 8'b00100000;
		color_arr[5697] = 8'b00100000;
		color_arr[5698] = 8'b00100000;
		color_arr[5699] = 8'b00100000;
		color_arr[5700] = 8'b00100000;
		color_arr[5701] = 8'b00100000;
		color_arr[5702] = 8'b00100000;
		color_arr[5703] = 8'b00100000;
		color_arr[5704] = 8'b00100000;
		color_arr[5705] = 8'b00100000;
		color_arr[5706] = 8'b00100000;
		color_arr[5707] = 8'b00100000;
		color_arr[5708] = 8'b00100000;
		color_arr[5709] = 8'b00100000;
		color_arr[5710] = 8'b00100000;
		color_arr[5711] = 8'b00100000;
		color_arr[5712] = 8'b00001000;
		color_arr[5713] = 8'b00001000;
		color_arr[5714] = 8'b00001000;
		color_arr[5715] = 8'b00001000;
		color_arr[5716] = 8'b00001000;
		color_arr[5717] = 8'b00001000;
		color_arr[5718] = 8'b00001000;
		color_arr[5719] = 8'b00001000;
		color_arr[5720] = 8'b00001000;
		color_arr[5721] = 8'b00001000;
		color_arr[5722] = 8'b00001000;
		color_arr[5723] = 8'b00001000;
		color_arr[5724] = 8'b00001000;
		color_arr[5725] = 8'b00001000;
		color_arr[5726] = 8'b00001000;
		color_arr[5727] = 8'b00001000;
		color_arr[5728] = 8'b00001000;
		color_arr[5729] = 8'b00000000;
		color_arr[5730] = 8'b00000000;
		color_arr[5731] = 8'b00000000;
		color_arr[5732] = 8'b00000000;
		color_arr[5733] = 8'b00001000;
		color_arr[5734] = 8'b00001000;
		color_arr[5735] = 8'b00001000;
		color_arr[5736] = 8'b00001000;
		color_arr[5737] = 8'b00001000;
		color_arr[5738] = 8'b00001000;
		color_arr[5739] = 8'b00001000;
		color_arr[5740] = 8'b00001000;
		color_arr[5741] = 8'b00001000;
		color_arr[5742] = 8'b00001000;
		color_arr[5743] = 8'b00001000;
		color_arr[5744] = 8'b00001000;
		color_arr[5745] = 8'b00001000;
		color_arr[5746] = 8'b00001000;
		color_arr[5747] = 8'b00001000;
		color_arr[5748] = 8'b00000000;
		color_arr[5749] = 8'b00000000;
		color_arr[5750] = 8'b00000000;
		color_arr[5751] = 8'b00001000;
		color_arr[5752] = 8'b00001000;
		color_arr[5753] = 8'b00001000;
		color_arr[5754] = 8'b00001000;
		color_arr[5755] = 8'b00001000;
		color_arr[5756] = 8'b00001000;
		color_arr[5757] = 8'b00010010;
		color_arr[5758] = 8'b00010010;
		color_arr[5759] = 8'b00010010;
		color_arr[5760] = 8'b00010010;
		color_arr[5761] = 8'b00010010;
		color_arr[5762] = 8'b00000000;
		color_arr[5763] = 8'b00000000;
		color_arr[5764] = 8'b00010010;
		color_arr[5765] = 8'b00010010;
		color_arr[5766] = 8'b00010010;
		color_arr[5767] = 8'b00010010;
		color_arr[5768] = 8'b00000010;
		color_arr[5769] = 8'b00000010;
		color_arr[5770] = 8'b00000010;
		color_arr[5771] = 8'b00000010;
		color_arr[5772] = 8'b00000010;
		color_arr[5773] = 8'b00000010;
		color_arr[5774] = 8'b00000010;
		color_arr[5775] = 8'b00000010;
		color_arr[5776] = 8'b00000010;
		color_arr[5777] = 8'b00000010;
		color_arr[5778] = 8'b00000010;
		color_arr[5779] = 8'b00000010;
		color_arr[5780] = 8'b00000010;
		color_arr[5781] = 8'b00000010;
		color_arr[5782] = 8'b00000010;
		color_arr[5783] = 8'b00000010;
		color_arr[5784] = 8'b00000010;
		color_arr[5785] = 8'b00000000;
		color_arr[5786] = 8'b00000000;
		color_arr[5787] = 8'b00000010;
		color_arr[5788] = 8'b00000010;
		color_arr[5789] = 8'b00000010;
		color_arr[5790] = 8'b00000010;
		color_arr[5791] = 8'b00000010;
		color_arr[5792] = 8'b00000010;
		color_arr[5793] = 8'b00000010;
		color_arr[5794] = 8'b00000010;
		color_arr[5795] = 8'b00000010;
		color_arr[5796] = 8'b00000010;
		color_arr[5797] = 8'b00000010;
		color_arr[5798] = 8'b00100000;
		color_arr[5799] = 8'b00100000;
		color_arr[5800] = 8'b00100000;
		color_arr[5801] = 8'b00100000;
		color_arr[5802] = 8'b00100000;
		color_arr[5803] = 8'b00100000;
		color_arr[5804] = 8'b00100000;
		color_arr[5805] = 8'b00100000;
		color_arr[5806] = 8'b00100000;
		color_arr[5807] = 8'b00100000;
		color_arr[5808] = 8'b00100000;
		color_arr[5809] = 8'b00100000;
		color_arr[5810] = 8'b00100000;
		color_arr[5811] = 8'b00100000;
		color_arr[5812] = 8'b00100000;
		color_arr[5813] = 8'b00100000;
		color_arr[5814] = 8'b00100000;
		color_arr[5815] = 8'b00100000;
		color_arr[5816] = 8'b00100000;
		color_arr[5817] = 8'b00100000;
		color_arr[5818] = 8'b00100000;
		color_arr[5819] = 8'b00100000;
		color_arr[5820] = 8'b00100000;
		color_arr[5821] = 8'b00100000;
		color_arr[5822] = 8'b00100000;
		color_arr[5823] = 8'b00100000;
		color_arr[5824] = 8'b00100000;
		color_arr[5825] = 8'b00100000;
		color_arr[5826] = 8'b00100000;
		color_arr[5827] = 8'b00100000;
		color_arr[5828] = 8'b00100000;
		color_arr[5829] = 8'b00100000;
		color_arr[5830] = 8'b00100000;
		color_arr[5831] = 8'b00100000;
		color_arr[5832] = 8'b00100000;
		color_arr[5833] = 8'b00100000;
		color_arr[5834] = 8'b00100000;
		color_arr[5835] = 8'b00100000;
		color_arr[5836] = 8'b00100000;
		color_arr[5837] = 8'b00100000;
		color_arr[5838] = 8'b00100000;
		color_arr[5839] = 8'b00100000;
		color_arr[5840] = 8'b00001000;
		color_arr[5841] = 8'b00001000;
		color_arr[5842] = 8'b00001000;
		color_arr[5843] = 8'b00001000;
		color_arr[5844] = 8'b00001000;
		color_arr[5845] = 8'b00001000;
		color_arr[5846] = 8'b00001000;
		color_arr[5847] = 8'b00001000;
		color_arr[5848] = 8'b00001000;
		color_arr[5849] = 8'b00001000;
		color_arr[5850] = 8'b00001000;
		color_arr[5851] = 8'b00001000;
		color_arr[5852] = 8'b00001000;
		color_arr[5853] = 8'b00001000;
		color_arr[5854] = 8'b00001000;
		color_arr[5855] = 8'b00001000;
		color_arr[5856] = 8'b00001000;
		color_arr[5857] = 8'b00000000;
		color_arr[5858] = 8'b00000000;
		color_arr[5859] = 8'b00000000;
		color_arr[5860] = 8'b00000000;
		color_arr[5861] = 8'b00001000;
		color_arr[5862] = 8'b00001000;
		color_arr[5863] = 8'b00001000;
		color_arr[5864] = 8'b00001000;
		color_arr[5865] = 8'b00001000;
		color_arr[5866] = 8'b00001000;
		color_arr[5867] = 8'b00001000;
		color_arr[5868] = 8'b00001000;
		color_arr[5869] = 8'b00001000;
		color_arr[5870] = 8'b00001000;
		color_arr[5871] = 8'b00001000;
		color_arr[5872] = 8'b00001000;
		color_arr[5873] = 8'b00001000;
		color_arr[5874] = 8'b00001000;
		color_arr[5875] = 8'b00001000;
		color_arr[5876] = 8'b00000000;
		color_arr[5877] = 8'b00000000;
		color_arr[5878] = 8'b00001000;
		color_arr[5879] = 8'b00001000;
		color_arr[5880] = 8'b00001000;
		color_arr[5881] = 8'b00001000;
		color_arr[5882] = 8'b00001000;
		color_arr[5883] = 8'b00001000;
		color_arr[5884] = 8'b00001000;
		color_arr[5885] = 8'b00010010;
		color_arr[5886] = 8'b00010010;
		color_arr[5887] = 8'b00010010;
		color_arr[5888] = 8'b00010010;
		color_arr[5889] = 8'b00010010;
		color_arr[5890] = 8'b00000000;
		color_arr[5891] = 8'b00000000;
		color_arr[5892] = 8'b00010010;
		color_arr[5893] = 8'b00010010;
		color_arr[5894] = 8'b00010010;
		color_arr[5895] = 8'b00010010;
		color_arr[5896] = 8'b00000010;
		color_arr[5897] = 8'b00000010;
		color_arr[5898] = 8'b00000010;
		color_arr[5899] = 8'b00000010;
		color_arr[5900] = 8'b00000010;
		color_arr[5901] = 8'b00000010;
		color_arr[5902] = 8'b00000010;
		color_arr[5903] = 8'b00000010;
		color_arr[5904] = 8'b00000010;
		color_arr[5905] = 8'b00000010;
		color_arr[5906] = 8'b00000010;
		color_arr[5907] = 8'b00000010;
		color_arr[5908] = 8'b00000010;
		color_arr[5909] = 8'b00000010;
		color_arr[5910] = 8'b00000010;
		color_arr[5911] = 8'b00000010;
		color_arr[5912] = 8'b00000000;
		color_arr[5913] = 8'b00000000;
		color_arr[5914] = 8'b00000000;
		color_arr[5915] = 8'b00000010;
		color_arr[5916] = 8'b00000010;
		color_arr[5917] = 8'b00000010;
		color_arr[5918] = 8'b00000010;
		color_arr[5919] = 8'b00000010;
		color_arr[5920] = 8'b00000010;
		color_arr[5921] = 8'b00000010;
		color_arr[5922] = 8'b00000010;
		color_arr[5923] = 8'b00000010;
		color_arr[5924] = 8'b00000010;
		color_arr[5925] = 8'b00000010;
		color_arr[5926] = 8'b00100000;
		color_arr[5927] = 8'b00100000;
		color_arr[5928] = 8'b00100000;
		color_arr[5929] = 8'b00100000;
		color_arr[5930] = 8'b00100000;
		color_arr[5931] = 8'b00100000;
		color_arr[5932] = 8'b00100000;
		color_arr[5933] = 8'b00100000;
		color_arr[5934] = 8'b00100000;
		color_arr[5935] = 8'b00100000;
		color_arr[5936] = 8'b00100000;
		color_arr[5937] = 8'b00100000;
		color_arr[5938] = 8'b00100000;
		color_arr[5939] = 8'b00100000;
		color_arr[5940] = 8'b00100000;
		color_arr[5941] = 8'b00100000;
		color_arr[5942] = 8'b00100000;
		color_arr[5943] = 8'b00100000;
		color_arr[5944] = 8'b00100000;
		color_arr[5945] = 8'b00100000;
		color_arr[5946] = 8'b00100000;
		color_arr[5947] = 8'b00100000;
		color_arr[5948] = 8'b00100000;
		color_arr[5949] = 8'b00100000;
		color_arr[5950] = 8'b00100000;
		color_arr[5951] = 8'b00100000;
		color_arr[5952] = 8'b00100000;
		color_arr[5953] = 8'b00100000;
		color_arr[5954] = 8'b00100000;
		color_arr[5955] = 8'b00100000;
		color_arr[5956] = 8'b00100000;
		color_arr[5957] = 8'b00100000;
		color_arr[5958] = 8'b00100000;
		color_arr[5959] = 8'b00100000;
		color_arr[5960] = 8'b00100000;
		color_arr[5961] = 8'b00100000;
		color_arr[5962] = 8'b00100000;
		color_arr[5963] = 8'b00100000;
		color_arr[5964] = 8'b00100000;
		color_arr[5965] = 8'b00100000;
		color_arr[5966] = 8'b00100000;
		color_arr[5967] = 8'b00100000;
		color_arr[5968] = 8'b00001000;
		color_arr[5969] = 8'b00001000;
		color_arr[5970] = 8'b00001000;
		color_arr[5971] = 8'b00001000;
		color_arr[5972] = 8'b00001000;
		color_arr[5973] = 8'b00001000;
		color_arr[5974] = 8'b00001000;
		color_arr[5975] = 8'b00001000;
		color_arr[5976] = 8'b00001000;
		color_arr[5977] = 8'b00001000;
		color_arr[5978] = 8'b00001000;
		color_arr[5979] = 8'b00001000;
		color_arr[5980] = 8'b00001000;
		color_arr[5981] = 8'b00001000;
		color_arr[5982] = 8'b00001000;
		color_arr[5983] = 8'b00001000;
		color_arr[5984] = 8'b00001000;
		color_arr[5985] = 8'b00001000;
		color_arr[5986] = 8'b00000000;
		color_arr[5987] = 8'b00000000;
		color_arr[5988] = 8'b00000000;
		color_arr[5989] = 8'b00000000;
		color_arr[5990] = 8'b00001000;
		color_arr[5991] = 8'b00001000;
		color_arr[5992] = 8'b00001000;
		color_arr[5993] = 8'b00001000;
		color_arr[5994] = 8'b00001000;
		color_arr[5995] = 8'b00001000;
		color_arr[5996] = 8'b00001000;
		color_arr[5997] = 8'b00001000;
		color_arr[5998] = 8'b00001000;
		color_arr[5999] = 8'b00001000;
		color_arr[6000] = 8'b00001000;
		color_arr[6001] = 8'b00001000;
		color_arr[6002] = 8'b00001000;
		color_arr[6003] = 8'b00001000;
		color_arr[6004] = 8'b00000000;
		color_arr[6005] = 8'b00000000;
		color_arr[6006] = 8'b00001000;
		color_arr[6007] = 8'b00001000;
		color_arr[6008] = 8'b00001000;
		color_arr[6009] = 8'b00001000;
		color_arr[6010] = 8'b00001000;
		color_arr[6011] = 8'b00001000;
		color_arr[6012] = 8'b00001000;
		color_arr[6013] = 8'b00010010;
		color_arr[6014] = 8'b00010010;
		color_arr[6015] = 8'b00010010;
		color_arr[6016] = 8'b00010010;
		color_arr[6017] = 8'b00010010;
		color_arr[6018] = 8'b00000000;
		color_arr[6019] = 8'b00000000;
		color_arr[6020] = 8'b00010010;
		color_arr[6021] = 8'b00010010;
		color_arr[6022] = 8'b00010010;
		color_arr[6023] = 8'b00010010;
		color_arr[6024] = 8'b00000010;
		color_arr[6025] = 8'b00000010;
		color_arr[6026] = 8'b00000010;
		color_arr[6027] = 8'b00000010;
		color_arr[6028] = 8'b00000010;
		color_arr[6029] = 8'b00000010;
		color_arr[6030] = 8'b00000010;
		color_arr[6031] = 8'b00000010;
		color_arr[6032] = 8'b00000010;
		color_arr[6033] = 8'b00000010;
		color_arr[6034] = 8'b00000010;
		color_arr[6035] = 8'b00000010;
		color_arr[6036] = 8'b00000010;
		color_arr[6037] = 8'b00000010;
		color_arr[6038] = 8'b00000010;
		color_arr[6039] = 8'b00000010;
		color_arr[6040] = 8'b00000000;
		color_arr[6041] = 8'b00000000;
		color_arr[6042] = 8'b00000010;
		color_arr[6043] = 8'b00000010;
		color_arr[6044] = 8'b00000010;
		color_arr[6045] = 8'b00000010;
		color_arr[6046] = 8'b00000010;
		color_arr[6047] = 8'b00000010;
		color_arr[6048] = 8'b00000010;
		color_arr[6049] = 8'b00000010;
		color_arr[6050] = 8'b00000010;
		color_arr[6051] = 8'b00000010;
		color_arr[6052] = 8'b00000010;
		color_arr[6053] = 8'b00000010;
		color_arr[6054] = 8'b00100000;
		color_arr[6055] = 8'b00100000;
		color_arr[6056] = 8'b00100000;
		color_arr[6057] = 8'b00100000;
		color_arr[6058] = 8'b00100000;
		color_arr[6059] = 8'b00100000;
		color_arr[6060] = 8'b00100000;
		color_arr[6061] = 8'b00100000;
		color_arr[6062] = 8'b00100000;
		color_arr[6063] = 8'b00100000;
		color_arr[6064] = 8'b00100000;
		color_arr[6065] = 8'b00100000;
		color_arr[6066] = 8'b00100000;
		color_arr[6067] = 8'b00100000;
		color_arr[6068] = 8'b00100000;
		color_arr[6069] = 8'b00100000;
		color_arr[6070] = 8'b00100000;
		color_arr[6071] = 8'b00100000;
		color_arr[6072] = 8'b00100000;
		color_arr[6073] = 8'b00100000;
		color_arr[6074] = 8'b00100000;
		color_arr[6075] = 8'b00100000;
		color_arr[6076] = 8'b00100000;
		color_arr[6077] = 8'b00100000;
		color_arr[6078] = 8'b00100000;
		color_arr[6079] = 8'b00100000;
		color_arr[6080] = 8'b00100000;
		color_arr[6081] = 8'b00100000;
		color_arr[6082] = 8'b00100000;
		color_arr[6083] = 8'b00100000;
		color_arr[6084] = 8'b00100000;
		color_arr[6085] = 8'b00100000;
		color_arr[6086] = 8'b00100000;
		color_arr[6087] = 8'b00100000;
		color_arr[6088] = 8'b00100000;
		color_arr[6089] = 8'b00100000;
		color_arr[6090] = 8'b00100000;
		color_arr[6091] = 8'b00100000;
		color_arr[6092] = 8'b00100000;
		color_arr[6093] = 8'b00100000;
		color_arr[6094] = 8'b00100000;
		color_arr[6095] = 8'b00100000;
		color_arr[6096] = 8'b00001000;
		color_arr[6097] = 8'b00001000;
		color_arr[6098] = 8'b00001000;
		color_arr[6099] = 8'b00001000;
		color_arr[6100] = 8'b00001000;
		color_arr[6101] = 8'b00001000;
		color_arr[6102] = 8'b00001000;
		color_arr[6103] = 8'b00001000;
		color_arr[6104] = 8'b00001000;
		color_arr[6105] = 8'b00001000;
		color_arr[6106] = 8'b00001000;
		color_arr[6107] = 8'b00001000;
		color_arr[6108] = 8'b00001000;
		color_arr[6109] = 8'b00001000;
		color_arr[6110] = 8'b00001000;
		color_arr[6111] = 8'b00001000;
		color_arr[6112] = 8'b00001000;
		color_arr[6113] = 8'b00001000;
		color_arr[6114] = 8'b00000000;
		color_arr[6115] = 8'b00000000;
		color_arr[6116] = 8'b00000000;
		color_arr[6117] = 8'b00000000;
		color_arr[6118] = 8'b00000000;
		color_arr[6119] = 8'b00001000;
		color_arr[6120] = 8'b00001000;
		color_arr[6121] = 8'b00001000;
		color_arr[6122] = 8'b00001000;
		color_arr[6123] = 8'b00001000;
		color_arr[6124] = 8'b00001000;
		color_arr[6125] = 8'b00001000;
		color_arr[6126] = 8'b00001000;
		color_arr[6127] = 8'b00001000;
		color_arr[6128] = 8'b00001000;
		color_arr[6129] = 8'b00001000;
		color_arr[6130] = 8'b00001000;
		color_arr[6131] = 8'b00001000;
		color_arr[6132] = 8'b00000000;
		color_arr[6133] = 8'b00000000;
		color_arr[6134] = 8'b00001000;
		color_arr[6135] = 8'b00001000;
		color_arr[6136] = 8'b00001000;
		color_arr[6137] = 8'b00001000;
		color_arr[6138] = 8'b00001000;
		color_arr[6139] = 8'b00001000;
		color_arr[6140] = 8'b00001000;
		color_arr[6141] = 8'b00010010;
		color_arr[6142] = 8'b00010010;
		color_arr[6143] = 8'b00010010;
		color_arr[6144] = 8'b00010010;
		color_arr[6145] = 8'b00010010;
		color_arr[6146] = 8'b00000000;
		color_arr[6147] = 8'b00000000;
		color_arr[6148] = 8'b00010010;
		color_arr[6149] = 8'b00010010;
		color_arr[6150] = 8'b00010010;
		color_arr[6151] = 8'b00010010;
		color_arr[6152] = 8'b00000010;
		color_arr[6153] = 8'b00000010;
		color_arr[6154] = 8'b00000010;
		color_arr[6155] = 8'b00000010;
		color_arr[6156] = 8'b00000010;
		color_arr[6157] = 8'b00000010;
		color_arr[6158] = 8'b00000010;
		color_arr[6159] = 8'b00000010;
		color_arr[6160] = 8'b00000010;
		color_arr[6161] = 8'b00000010;
		color_arr[6162] = 8'b00000010;
		color_arr[6163] = 8'b00000010;
		color_arr[6164] = 8'b00000010;
		color_arr[6165] = 8'b00000010;
		color_arr[6166] = 8'b00000010;
		color_arr[6167] = 8'b00000000;
		color_arr[6168] = 8'b00000000;
		color_arr[6169] = 8'b00000000;
		color_arr[6170] = 8'b00000010;
		color_arr[6171] = 8'b00000010;
		color_arr[6172] = 8'b00000010;
		color_arr[6173] = 8'b00000010;
		color_arr[6174] = 8'b00000010;
		color_arr[6175] = 8'b00000010;
		color_arr[6176] = 8'b00000010;
		color_arr[6177] = 8'b00000010;
		color_arr[6178] = 8'b00000010;
		color_arr[6179] = 8'b00000010;
		color_arr[6180] = 8'b00000010;
		color_arr[6181] = 8'b00000010;
		color_arr[6182] = 8'b00100000;
		color_arr[6183] = 8'b00100000;
		color_arr[6184] = 8'b00100000;
		color_arr[6185] = 8'b00100000;
		color_arr[6186] = 8'b00100000;
		color_arr[6187] = 8'b00100000;
		color_arr[6188] = 8'b00100000;
		color_arr[6189] = 8'b00100000;
		color_arr[6190] = 8'b00100000;
		color_arr[6191] = 8'b00100000;
		color_arr[6192] = 8'b00100000;
		color_arr[6193] = 8'b00100000;
		color_arr[6194] = 8'b00100000;
		color_arr[6195] = 8'b00100000;
		color_arr[6196] = 8'b00100000;
		color_arr[6197] = 8'b00100000;
		color_arr[6198] = 8'b00100000;
		color_arr[6199] = 8'b00100000;
		color_arr[6200] = 8'b00100000;
		color_arr[6201] = 8'b00100000;
		color_arr[6202] = 8'b00100000;
		color_arr[6203] = 8'b00100000;
		color_arr[6204] = 8'b00100000;
		color_arr[6205] = 8'b00100000;
		color_arr[6206] = 8'b00100000;
		color_arr[6207] = 8'b00100000;
		color_arr[6208] = 8'b00100000;
		color_arr[6209] = 8'b00100000;
		color_arr[6210] = 8'b00100000;
		color_arr[6211] = 8'b00100000;
		color_arr[6212] = 8'b00100000;
		color_arr[6213] = 8'b00100000;
		color_arr[6214] = 8'b00100000;
		color_arr[6215] = 8'b00100000;
		color_arr[6216] = 8'b00100000;
		color_arr[6217] = 8'b00100000;
		color_arr[6218] = 8'b00100000;
		color_arr[6219] = 8'b00100000;
		color_arr[6220] = 8'b00100000;
		color_arr[6221] = 8'b00100000;
		color_arr[6222] = 8'b00100000;
		color_arr[6223] = 8'b00100000;
		color_arr[6224] = 8'b00001000;
		color_arr[6225] = 8'b00001000;
		color_arr[6226] = 8'b00001000;
		color_arr[6227] = 8'b00001000;
		color_arr[6228] = 8'b00001000;
		color_arr[6229] = 8'b00001000;
		color_arr[6230] = 8'b00001000;
		color_arr[6231] = 8'b00001000;
		color_arr[6232] = 8'b00001000;
		color_arr[6233] = 8'b00001000;
		color_arr[6234] = 8'b00001000;
		color_arr[6235] = 8'b00001000;
		color_arr[6236] = 8'b00001000;
		color_arr[6237] = 8'b00001000;
		color_arr[6238] = 8'b00001000;
		color_arr[6239] = 8'b00001000;
		color_arr[6240] = 8'b00001000;
		color_arr[6241] = 8'b00001000;
		color_arr[6242] = 8'b00000000;
		color_arr[6243] = 8'b00000000;
		color_arr[6244] = 8'b00001000;
		color_arr[6245] = 8'b00000000;
		color_arr[6246] = 8'b00000000;
		color_arr[6247] = 8'b00000000;
		color_arr[6248] = 8'b00001000;
		color_arr[6249] = 8'b00001000;
		color_arr[6250] = 8'b00001000;
		color_arr[6251] = 8'b00001000;
		color_arr[6252] = 8'b00001000;
		color_arr[6253] = 8'b00001000;
		color_arr[6254] = 8'b00001000;
		color_arr[6255] = 8'b00001000;
		color_arr[6256] = 8'b00001000;
		color_arr[6257] = 8'b00001000;
		color_arr[6258] = 8'b00001000;
		color_arr[6259] = 8'b00001000;
		color_arr[6260] = 8'b00000000;
		color_arr[6261] = 8'b00000000;
		color_arr[6262] = 8'b00001000;
		color_arr[6263] = 8'b00001000;
		color_arr[6264] = 8'b00001000;
		color_arr[6265] = 8'b00001000;
		color_arr[6266] = 8'b00001000;
		color_arr[6267] = 8'b00001000;
		color_arr[6268] = 8'b00001000;
		color_arr[6269] = 8'b00010010;
		color_arr[6270] = 8'b00010010;
		color_arr[6271] = 8'b00010010;
		color_arr[6272] = 8'b00010010;
		color_arr[6273] = 8'b00010010;
		color_arr[6274] = 8'b00000000;
		color_arr[6275] = 8'b00000000;
		color_arr[6276] = 8'b00010010;
		color_arr[6277] = 8'b00010010;
		color_arr[6278] = 8'b00010010;
		color_arr[6279] = 8'b00010010;
		color_arr[6280] = 8'b00000010;
		color_arr[6281] = 8'b00000010;
		color_arr[6282] = 8'b00000010;
		color_arr[6283] = 8'b00000010;
		color_arr[6284] = 8'b00000010;
		color_arr[6285] = 8'b00000010;
		color_arr[6286] = 8'b00000010;
		color_arr[6287] = 8'b00000010;
		color_arr[6288] = 8'b00000010;
		color_arr[6289] = 8'b00000010;
		color_arr[6290] = 8'b00000010;
		color_arr[6291] = 8'b00000010;
		color_arr[6292] = 8'b00000010;
		color_arr[6293] = 8'b00000010;
		color_arr[6294] = 8'b00000010;
		color_arr[6295] = 8'b00000000;
		color_arr[6296] = 8'b00000000;
		color_arr[6297] = 8'b00000010;
		color_arr[6298] = 8'b00000010;
		color_arr[6299] = 8'b00000010;
		color_arr[6300] = 8'b00000010;
		color_arr[6301] = 8'b00000010;
		color_arr[6302] = 8'b00000010;
		color_arr[6303] = 8'b00000010;
		color_arr[6304] = 8'b00000010;
		color_arr[6305] = 8'b00000010;
		color_arr[6306] = 8'b00000010;
		color_arr[6307] = 8'b00000010;
		color_arr[6308] = 8'b00000010;
		color_arr[6309] = 8'b00000010;
		color_arr[6310] = 8'b00100000;
		color_arr[6311] = 8'b00100000;
		color_arr[6312] = 8'b00100000;
		color_arr[6313] = 8'b00100000;
		color_arr[6314] = 8'b00100000;
		color_arr[6315] = 8'b00100000;
		color_arr[6316] = 8'b00100000;
		color_arr[6317] = 8'b00100000;
		color_arr[6318] = 8'b00100000;
		color_arr[6319] = 8'b00100000;
		color_arr[6320] = 8'b00100000;
		color_arr[6321] = 8'b00100000;
		color_arr[6322] = 8'b00100000;
		color_arr[6323] = 8'b00100000;
		color_arr[6324] = 8'b00100000;
		color_arr[6325] = 8'b00100000;
		color_arr[6326] = 8'b00100000;
		color_arr[6327] = 8'b00100000;
		color_arr[6328] = 8'b00100000;
		color_arr[6329] = 8'b00100000;
		color_arr[6330] = 8'b00100000;
		color_arr[6331] = 8'b00100000;
		color_arr[6332] = 8'b00100000;
		color_arr[6333] = 8'b00100000;
		color_arr[6334] = 8'b00100000;
		color_arr[6335] = 8'b00100000;
		color_arr[6336] = 8'b00100000;
		color_arr[6337] = 8'b00100000;
		color_arr[6338] = 8'b00100000;
		color_arr[6339] = 8'b00100000;
		color_arr[6340] = 8'b00100000;
		color_arr[6341] = 8'b00100000;
		color_arr[6342] = 8'b00100000;
		color_arr[6343] = 8'b00100000;
		color_arr[6344] = 8'b00100000;
		color_arr[6345] = 8'b00100000;
		color_arr[6346] = 8'b00100000;
		color_arr[6347] = 8'b00100000;
		color_arr[6348] = 8'b00100000;
		color_arr[6349] = 8'b00100000;
		color_arr[6350] = 8'b00100000;
		color_arr[6351] = 8'b00100000;
		color_arr[6352] = 8'b00001000;
		color_arr[6353] = 8'b00001000;
		color_arr[6354] = 8'b00001000;
		color_arr[6355] = 8'b00001000;
		color_arr[6356] = 8'b00001000;
		color_arr[6357] = 8'b00001000;
		color_arr[6358] = 8'b00001000;
		color_arr[6359] = 8'b00001000;
		color_arr[6360] = 8'b00001000;
		color_arr[6361] = 8'b00001000;
		color_arr[6362] = 8'b00001000;
		color_arr[6363] = 8'b00001000;
		color_arr[6364] = 8'b00001000;
		color_arr[6365] = 8'b00001000;
		color_arr[6366] = 8'b00001000;
		color_arr[6367] = 8'b00001000;
		color_arr[6368] = 8'b00001000;
		color_arr[6369] = 8'b00001000;
		color_arr[6370] = 8'b00000000;
		color_arr[6371] = 8'b00000000;
		color_arr[6372] = 8'b00001000;
		color_arr[6373] = 8'b00001000;
		color_arr[6374] = 8'b00000000;
		color_arr[6375] = 8'b00000000;
		color_arr[6376] = 8'b00000000;
		color_arr[6377] = 8'b00000000;
		color_arr[6378] = 8'b00001000;
		color_arr[6379] = 8'b00001000;
		color_arr[6380] = 8'b00001000;
		color_arr[6381] = 8'b00001000;
		color_arr[6382] = 8'b00001000;
		color_arr[6383] = 8'b00001000;
		color_arr[6384] = 8'b00001000;
		color_arr[6385] = 8'b00001000;
		color_arr[6386] = 8'b00001000;
		color_arr[6387] = 8'b00001000;
		color_arr[6388] = 8'b00000000;
		color_arr[6389] = 8'b00000000;
		color_arr[6390] = 8'b00001000;
		color_arr[6391] = 8'b00001000;
		color_arr[6392] = 8'b00001000;
		color_arr[6393] = 8'b00001000;
		color_arr[6394] = 8'b00001000;
		color_arr[6395] = 8'b00001000;
		color_arr[6396] = 8'b00001000;
		color_arr[6397] = 8'b00010010;
		color_arr[6398] = 8'b00010010;
		color_arr[6399] = 8'b00010010;
		color_arr[6400] = 8'b00010010;
		color_arr[6401] = 8'b00010010;
		color_arr[6402] = 8'b00000000;
		color_arr[6403] = 8'b00000000;
		color_arr[6404] = 8'b00010010;
		color_arr[6405] = 8'b00010010;
		color_arr[6406] = 8'b00010010;
		color_arr[6407] = 8'b00010010;
		color_arr[6408] = 8'b00000010;
		color_arr[6409] = 8'b00000010;
		color_arr[6410] = 8'b00000010;
		color_arr[6411] = 8'b00000010;
		color_arr[6412] = 8'b00000010;
		color_arr[6413] = 8'b00000010;
		color_arr[6414] = 8'b00000010;
		color_arr[6415] = 8'b00000010;
		color_arr[6416] = 8'b00000010;
		color_arr[6417] = 8'b00000010;
		color_arr[6418] = 8'b00000010;
		color_arr[6419] = 8'b00000010;
		color_arr[6420] = 8'b00000010;
		color_arr[6421] = 8'b00000010;
		color_arr[6422] = 8'b00000000;
		color_arr[6423] = 8'b00000000;
		color_arr[6424] = 8'b00000000;
		color_arr[6425] = 8'b00000010;
		color_arr[6426] = 8'b00000010;
		color_arr[6427] = 8'b00000010;
		color_arr[6428] = 8'b00000010;
		color_arr[6429] = 8'b00000010;
		color_arr[6430] = 8'b00000010;
		color_arr[6431] = 8'b00000010;
		color_arr[6432] = 8'b00000010;
		color_arr[6433] = 8'b00000010;
		color_arr[6434] = 8'b00000010;
		color_arr[6435] = 8'b00000010;
		color_arr[6436] = 8'b00000010;
		color_arr[6437] = 8'b00000010;
		color_arr[6438] = 8'b00100000;
		color_arr[6439] = 8'b00100000;
		color_arr[6440] = 8'b00100000;
		color_arr[6441] = 8'b00100000;
		color_arr[6442] = 8'b00100000;
		color_arr[6443] = 8'b00100000;
		color_arr[6444] = 8'b00100000;
		color_arr[6445] = 8'b00100000;
		color_arr[6446] = 8'b00100000;
		color_arr[6447] = 8'b00100000;
		color_arr[6448] = 8'b00100000;
		color_arr[6449] = 8'b00100000;
		color_arr[6450] = 8'b00100000;
		color_arr[6451] = 8'b00100000;
		color_arr[6452] = 8'b00100000;
		color_arr[6453] = 8'b00100000;
		color_arr[6454] = 8'b00100000;
		color_arr[6455] = 8'b00100000;
		color_arr[6456] = 8'b00100000;
		color_arr[6457] = 8'b00100000;
		color_arr[6458] = 8'b00100000;
		color_arr[6459] = 8'b00100000;
		color_arr[6460] = 8'b00100000;
		color_arr[6461] = 8'b00100000;
		color_arr[6462] = 8'b00100000;
		color_arr[6463] = 8'b00100000;
		color_arr[6464] = 8'b00100000;
		color_arr[6465] = 8'b00100000;
		color_arr[6466] = 8'b00100000;
		color_arr[6467] = 8'b00100000;
		color_arr[6468] = 8'b00100000;
		color_arr[6469] = 8'b00100000;
		color_arr[6470] = 8'b00100000;
		color_arr[6471] = 8'b00100000;
		color_arr[6472] = 8'b00100000;
		color_arr[6473] = 8'b00100000;
		color_arr[6474] = 8'b00100000;
		color_arr[6475] = 8'b00100000;
		color_arr[6476] = 8'b00100000;
		color_arr[6477] = 8'b00100000;
		color_arr[6478] = 8'b00100000;
		color_arr[6479] = 8'b00100000;
		color_arr[6480] = 8'b00001000;
		color_arr[6481] = 8'b00001000;
		color_arr[6482] = 8'b00001000;
		color_arr[6483] = 8'b00001000;
		color_arr[6484] = 8'b00001000;
		color_arr[6485] = 8'b00001000;
		color_arr[6486] = 8'b00001000;
		color_arr[6487] = 8'b00001000;
		color_arr[6488] = 8'b00001000;
		color_arr[6489] = 8'b00001000;
		color_arr[6490] = 8'b00001000;
		color_arr[6491] = 8'b00001000;
		color_arr[6492] = 8'b00001000;
		color_arr[6493] = 8'b00001000;
		color_arr[6494] = 8'b00001000;
		color_arr[6495] = 8'b00001000;
		color_arr[6496] = 8'b00001000;
		color_arr[6497] = 8'b00001000;
		color_arr[6498] = 8'b00000000;
		color_arr[6499] = 8'b00000000;
		color_arr[6500] = 8'b00001000;
		color_arr[6501] = 8'b00001000;
		color_arr[6502] = 8'b00001000;
		color_arr[6503] = 8'b00000000;
		color_arr[6504] = 8'b00000000;
		color_arr[6505] = 8'b00000000;
		color_arr[6506] = 8'b00000000;
		color_arr[6507] = 8'b00001000;
		color_arr[6508] = 8'b00001000;
		color_arr[6509] = 8'b00001000;
		color_arr[6510] = 8'b00001000;
		color_arr[6511] = 8'b00001000;
		color_arr[6512] = 8'b00001000;
		color_arr[6513] = 8'b00001000;
		color_arr[6514] = 8'b00001000;
		color_arr[6515] = 8'b00001000;
		color_arr[6516] = 8'b00000000;
		color_arr[6517] = 8'b00000000;
		color_arr[6518] = 8'b00001000;
		color_arr[6519] = 8'b00001000;
		color_arr[6520] = 8'b00001000;
		color_arr[6521] = 8'b00001000;
		color_arr[6522] = 8'b00001000;
		color_arr[6523] = 8'b00001000;
		color_arr[6524] = 8'b00001000;
		color_arr[6525] = 8'b00010010;
		color_arr[6526] = 8'b00010010;
		color_arr[6527] = 8'b00010010;
		color_arr[6528] = 8'b00010010;
		color_arr[6529] = 8'b00010010;
		color_arr[6530] = 8'b00000000;
		color_arr[6531] = 8'b00000000;
		color_arr[6532] = 8'b00010010;
		color_arr[6533] = 8'b00010010;
		color_arr[6534] = 8'b00010010;
		color_arr[6535] = 8'b00010010;
		color_arr[6536] = 8'b00000010;
		color_arr[6537] = 8'b00000010;
		color_arr[6538] = 8'b00000010;
		color_arr[6539] = 8'b00000010;
		color_arr[6540] = 8'b00000010;
		color_arr[6541] = 8'b00000010;
		color_arr[6542] = 8'b00000010;
		color_arr[6543] = 8'b00000010;
		color_arr[6544] = 8'b00000010;
		color_arr[6545] = 8'b00000010;
		color_arr[6546] = 8'b00000010;
		color_arr[6547] = 8'b00000010;
		color_arr[6548] = 8'b00000010;
		color_arr[6549] = 8'b00000010;
		color_arr[6550] = 8'b00000000;
		color_arr[6551] = 8'b00000000;
		color_arr[6552] = 8'b00000010;
		color_arr[6553] = 8'b00000010;
		color_arr[6554] = 8'b00000010;
		color_arr[6555] = 8'b00000010;
		color_arr[6556] = 8'b00000010;
		color_arr[6557] = 8'b00000010;
		color_arr[6558] = 8'b00000010;
		color_arr[6559] = 8'b00000010;
		color_arr[6560] = 8'b00000010;
		color_arr[6561] = 8'b00000010;
		color_arr[6562] = 8'b00000010;
		color_arr[6563] = 8'b00000010;
		color_arr[6564] = 8'b00000010;
		color_arr[6565] = 8'b00000010;
		color_arr[6566] = 8'b00100000;
		color_arr[6567] = 8'b00100000;
		color_arr[6568] = 8'b00100000;
		color_arr[6569] = 8'b00100000;
		color_arr[6570] = 8'b00100000;
		color_arr[6571] = 8'b00100000;
		color_arr[6572] = 8'b00100000;
		color_arr[6573] = 8'b00100000;
		color_arr[6574] = 8'b00100000;
		color_arr[6575] = 8'b00100000;
		color_arr[6576] = 8'b00100000;
		color_arr[6577] = 8'b00100000;
		color_arr[6578] = 8'b00100000;
		color_arr[6579] = 8'b00100000;
		color_arr[6580] = 8'b00100000;
		color_arr[6581] = 8'b00100000;
		color_arr[6582] = 8'b00100000;
		color_arr[6583] = 8'b00100000;
		color_arr[6584] = 8'b00100000;
		color_arr[6585] = 8'b00100000;
		color_arr[6586] = 8'b00100000;
		color_arr[6587] = 8'b00100000;
		color_arr[6588] = 8'b00100000;
		color_arr[6589] = 8'b00100000;
		color_arr[6590] = 8'b00100000;
		color_arr[6591] = 8'b00100000;
		color_arr[6592] = 8'b00100000;
		color_arr[6593] = 8'b00100000;
		color_arr[6594] = 8'b00100000;
		color_arr[6595] = 8'b00100000;
		color_arr[6596] = 8'b00100000;
		color_arr[6597] = 8'b00100000;
		color_arr[6598] = 8'b00100000;
		color_arr[6599] = 8'b00100000;
		color_arr[6600] = 8'b00100000;
		color_arr[6601] = 8'b00100000;
		color_arr[6602] = 8'b00100000;
		color_arr[6603] = 8'b00100000;
		color_arr[6604] = 8'b00100000;
		color_arr[6605] = 8'b00100000;
		color_arr[6606] = 8'b00100000;
		color_arr[6607] = 8'b00100000;
		color_arr[6608] = 8'b00001000;
		color_arr[6609] = 8'b00001000;
		color_arr[6610] = 8'b00001000;
		color_arr[6611] = 8'b00001000;
		color_arr[6612] = 8'b00001000;
		color_arr[6613] = 8'b00001000;
		color_arr[6614] = 8'b00001000;
		color_arr[6615] = 8'b00001000;
		color_arr[6616] = 8'b00001000;
		color_arr[6617] = 8'b00001000;
		color_arr[6618] = 8'b00001000;
		color_arr[6619] = 8'b00001000;
		color_arr[6620] = 8'b00001000;
		color_arr[6621] = 8'b00001000;
		color_arr[6622] = 8'b00001000;
		color_arr[6623] = 8'b00001000;
		color_arr[6624] = 8'b00001000;
		color_arr[6625] = 8'b00000000;
		color_arr[6626] = 8'b00000000;
		color_arr[6627] = 8'b00000000;
		color_arr[6628] = 8'b00001000;
		color_arr[6629] = 8'b00001000;
		color_arr[6630] = 8'b00001000;
		color_arr[6631] = 8'b00001000;
		color_arr[6632] = 8'b00001000;
		color_arr[6633] = 8'b00000000;
		color_arr[6634] = 8'b00000000;
		color_arr[6635] = 8'b00000000;
		color_arr[6636] = 8'b00001000;
		color_arr[6637] = 8'b00001000;
		color_arr[6638] = 8'b00001000;
		color_arr[6639] = 8'b00001000;
		color_arr[6640] = 8'b00001000;
		color_arr[6641] = 8'b00001000;
		color_arr[6642] = 8'b00001000;
		color_arr[6643] = 8'b00001000;
		color_arr[6644] = 8'b00000000;
		color_arr[6645] = 8'b00000000;
		color_arr[6646] = 8'b00001000;
		color_arr[6647] = 8'b00001000;
		color_arr[6648] = 8'b00001000;
		color_arr[6649] = 8'b00001000;
		color_arr[6650] = 8'b00001000;
		color_arr[6651] = 8'b00001000;
		color_arr[6652] = 8'b00001000;
		color_arr[6653] = 8'b00010010;
		color_arr[6654] = 8'b00010010;
		color_arr[6655] = 8'b00010010;
		color_arr[6656] = 8'b00010010;
		color_arr[6657] = 8'b00010010;
		color_arr[6658] = 8'b00000000;
		color_arr[6659] = 8'b00000000;
		color_arr[6660] = 8'b00010010;
		color_arr[6661] = 8'b00010010;
		color_arr[6662] = 8'b00010010;
		color_arr[6663] = 8'b00010010;
		color_arr[6664] = 8'b00000010;
		color_arr[6665] = 8'b00000010;
		color_arr[6666] = 8'b00000010;
		color_arr[6667] = 8'b00000010;
		color_arr[6668] = 8'b00000010;
		color_arr[6669] = 8'b00000010;
		color_arr[6670] = 8'b00000010;
		color_arr[6671] = 8'b00000010;
		color_arr[6672] = 8'b00000010;
		color_arr[6673] = 8'b00000010;
		color_arr[6674] = 8'b00000010;
		color_arr[6675] = 8'b00000010;
		color_arr[6676] = 8'b00000010;
		color_arr[6677] = 8'b00000010;
		color_arr[6678] = 8'b00000000;
		color_arr[6679] = 8'b00000000;
		color_arr[6680] = 8'b00000010;
		color_arr[6681] = 8'b00000010;
		color_arr[6682] = 8'b00000010;
		color_arr[6683] = 8'b00000010;
		color_arr[6684] = 8'b00000010;
		color_arr[6685] = 8'b00000010;
		color_arr[6686] = 8'b00000010;
		color_arr[6687] = 8'b00000010;
		color_arr[6688] = 8'b00000010;
		color_arr[6689] = 8'b00000010;
		color_arr[6690] = 8'b00000010;
		color_arr[6691] = 8'b00000010;
		color_arr[6692] = 8'b00000010;
		color_arr[6693] = 8'b00000010;
		color_arr[6694] = 8'b00100000;
		color_arr[6695] = 8'b00100000;
		color_arr[6696] = 8'b00100000;
		color_arr[6697] = 8'b00100000;
		color_arr[6698] = 8'b00100000;
		color_arr[6699] = 8'b00100000;
		color_arr[6700] = 8'b00100000;
		color_arr[6701] = 8'b00100000;
		color_arr[6702] = 8'b00100000;
		color_arr[6703] = 8'b00100000;
		color_arr[6704] = 8'b00100000;
		color_arr[6705] = 8'b00100000;
		color_arr[6706] = 8'b00100000;
		color_arr[6707] = 8'b00100000;
		color_arr[6708] = 8'b00100000;
		color_arr[6709] = 8'b00100000;
		color_arr[6710] = 8'b00100000;
		color_arr[6711] = 8'b00100000;
		color_arr[6712] = 8'b00100000;
		color_arr[6713] = 8'b00100000;
		color_arr[6714] = 8'b00100000;
		color_arr[6715] = 8'b00100000;
		color_arr[6716] = 8'b00100000;
		color_arr[6717] = 8'b00100000;
		color_arr[6718] = 8'b00100000;
		color_arr[6719] = 8'b00100000;
		color_arr[6720] = 8'b00100000;
		color_arr[6721] = 8'b00100000;
		color_arr[6722] = 8'b00100000;
		color_arr[6723] = 8'b00100000;
		color_arr[6724] = 8'b00100000;
		color_arr[6725] = 8'b00100000;
		color_arr[6726] = 8'b00100000;
		color_arr[6727] = 8'b00100000;
		color_arr[6728] = 8'b00100000;
		color_arr[6729] = 8'b00100000;
		color_arr[6730] = 8'b00100000;
		color_arr[6731] = 8'b00100000;
		color_arr[6732] = 8'b00100000;
		color_arr[6733] = 8'b00100000;
		color_arr[6734] = 8'b00100000;
		color_arr[6735] = 8'b00100000;
		color_arr[6736] = 8'b00001000;
		color_arr[6737] = 8'b00001000;
		color_arr[6738] = 8'b00001000;
		color_arr[6739] = 8'b00001000;
		color_arr[6740] = 8'b00001000;
		color_arr[6741] = 8'b00001000;
		color_arr[6742] = 8'b00001000;
		color_arr[6743] = 8'b00001000;
		color_arr[6744] = 8'b00001000;
		color_arr[6745] = 8'b00001000;
		color_arr[6746] = 8'b00001000;
		color_arr[6747] = 8'b00001000;
		color_arr[6748] = 8'b00001000;
		color_arr[6749] = 8'b00001000;
		color_arr[6750] = 8'b00001000;
		color_arr[6751] = 8'b00001000;
		color_arr[6752] = 8'b00001000;
		color_arr[6753] = 8'b00000000;
		color_arr[6754] = 8'b00000000;
		color_arr[6755] = 8'b00001000;
		color_arr[6756] = 8'b00001000;
		color_arr[6757] = 8'b00001000;
		color_arr[6758] = 8'b00001000;
		color_arr[6759] = 8'b00001000;
		color_arr[6760] = 8'b00001000;
		color_arr[6761] = 8'b00001000;
		color_arr[6762] = 8'b00000000;
		color_arr[6763] = 8'b00000000;
		color_arr[6764] = 8'b00000000;
		color_arr[6765] = 8'b00001000;
		color_arr[6766] = 8'b00001000;
		color_arr[6767] = 8'b00001000;
		color_arr[6768] = 8'b00001000;
		color_arr[6769] = 8'b00001000;
		color_arr[6770] = 8'b00001000;
		color_arr[6771] = 8'b00001000;
		color_arr[6772] = 8'b00000000;
		color_arr[6773] = 8'b00000000;
		color_arr[6774] = 8'b00001000;
		color_arr[6775] = 8'b00001000;
		color_arr[6776] = 8'b00001000;
		color_arr[6777] = 8'b00001000;
		color_arr[6778] = 8'b00001000;
		color_arr[6779] = 8'b00001000;
		color_arr[6780] = 8'b00001000;
		color_arr[6781] = 8'b00010010;
		color_arr[6782] = 8'b00010010;
		color_arr[6783] = 8'b00010010;
		color_arr[6784] = 8'b00010010;
		color_arr[6785] = 8'b00010010;
		color_arr[6786] = 8'b00000000;
		color_arr[6787] = 8'b00000000;
		color_arr[6788] = 8'b00010010;
		color_arr[6789] = 8'b00010010;
		color_arr[6790] = 8'b00010010;
		color_arr[6791] = 8'b00010010;
		color_arr[6792] = 8'b00000010;
		color_arr[6793] = 8'b00000010;
		color_arr[6794] = 8'b00000010;
		color_arr[6795] = 8'b00000010;
		color_arr[6796] = 8'b00000010;
		color_arr[6797] = 8'b00000010;
		color_arr[6798] = 8'b00000010;
		color_arr[6799] = 8'b00000010;
		color_arr[6800] = 8'b00000010;
		color_arr[6801] = 8'b00000010;
		color_arr[6802] = 8'b00000010;
		color_arr[6803] = 8'b00000010;
		color_arr[6804] = 8'b00000010;
		color_arr[6805] = 8'b00000010;
		color_arr[6806] = 8'b00000000;
		color_arr[6807] = 8'b00000000;
		color_arr[6808] = 8'b00000010;
		color_arr[6809] = 8'b00000010;
		color_arr[6810] = 8'b00000010;
		color_arr[6811] = 8'b00000010;
		color_arr[6812] = 8'b00000010;
		color_arr[6813] = 8'b00000010;
		color_arr[6814] = 8'b00000010;
		color_arr[6815] = 8'b00000010;
		color_arr[6816] = 8'b00000010;
		color_arr[6817] = 8'b00000010;
		color_arr[6818] = 8'b00000010;
		color_arr[6819] = 8'b00000010;
		color_arr[6820] = 8'b00000010;
		color_arr[6821] = 8'b00000010;
		color_arr[6822] = 8'b00100000;
		color_arr[6823] = 8'b00100000;
		color_arr[6824] = 8'b00100000;
		color_arr[6825] = 8'b00100000;
		color_arr[6826] = 8'b00100000;
		color_arr[6827] = 8'b00100000;
		color_arr[6828] = 8'b00100000;
		color_arr[6829] = 8'b00100000;
		color_arr[6830] = 8'b00100000;
		color_arr[6831] = 8'b00100000;
		color_arr[6832] = 8'b00100000;
		color_arr[6833] = 8'b00100000;
		color_arr[6834] = 8'b00100000;
		color_arr[6835] = 8'b00100000;
		color_arr[6836] = 8'b00100000;
		color_arr[6837] = 8'b00100000;
		color_arr[6838] = 8'b00100000;
		color_arr[6839] = 8'b00100000;
		color_arr[6840] = 8'b00100000;
		color_arr[6841] = 8'b00100000;
		color_arr[6842] = 8'b00100000;
		color_arr[6843] = 8'b00100000;
		color_arr[6844] = 8'b00100000;
		color_arr[6845] = 8'b00100000;
		color_arr[6846] = 8'b00100000;
		color_arr[6847] = 8'b00100000;
		color_arr[6848] = 8'b00100000;
		color_arr[6849] = 8'b00100000;
		color_arr[6850] = 8'b00100000;
		color_arr[6851] = 8'b00100000;
		color_arr[6852] = 8'b00100000;
		color_arr[6853] = 8'b00100000;
		color_arr[6854] = 8'b00100000;
		color_arr[6855] = 8'b00100000;
		color_arr[6856] = 8'b00100000;
		color_arr[6857] = 8'b00100000;
		color_arr[6858] = 8'b00100000;
		color_arr[6859] = 8'b00100000;
		color_arr[6860] = 8'b00100000;
		color_arr[6861] = 8'b00100000;
		color_arr[6862] = 8'b00100000;
		color_arr[6863] = 8'b00100000;
		color_arr[6864] = 8'b00001000;
		color_arr[6865] = 8'b00001000;
		color_arr[6866] = 8'b00001000;
		color_arr[6867] = 8'b00001000;
		color_arr[6868] = 8'b00001000;
		color_arr[6869] = 8'b00001000;
		color_arr[6870] = 8'b00001000;
		color_arr[6871] = 8'b00001000;
		color_arr[6872] = 8'b00001000;
		color_arr[6873] = 8'b00001000;
		color_arr[6874] = 8'b00001000;
		color_arr[6875] = 8'b00001000;
		color_arr[6876] = 8'b00001000;
		color_arr[6877] = 8'b00001000;
		color_arr[6878] = 8'b00001000;
		color_arr[6879] = 8'b00001000;
		color_arr[6880] = 8'b00000000;
		color_arr[6881] = 8'b00000000;
		color_arr[6882] = 8'b00000000;
		color_arr[6883] = 8'b00001000;
		color_arr[6884] = 8'b00001000;
		color_arr[6885] = 8'b00001000;
		color_arr[6886] = 8'b00001000;
		color_arr[6887] = 8'b00001000;
		color_arr[6888] = 8'b00001000;
		color_arr[6889] = 8'b00001000;
		color_arr[6890] = 8'b00001000;
		color_arr[6891] = 8'b00000000;
		color_arr[6892] = 8'b00000000;
		color_arr[6893] = 8'b00001000;
		color_arr[6894] = 8'b00001000;
		color_arr[6895] = 8'b00001000;
		color_arr[6896] = 8'b00001000;
		color_arr[6897] = 8'b00001000;
		color_arr[6898] = 8'b00001000;
		color_arr[6899] = 8'b00001000;
		color_arr[6900] = 8'b00000000;
		color_arr[6901] = 8'b00000000;
		color_arr[6902] = 8'b00001000;
		color_arr[6903] = 8'b00001000;
		color_arr[6904] = 8'b00001000;
		color_arr[6905] = 8'b00001000;
		color_arr[6906] = 8'b00001000;
		color_arr[6907] = 8'b00001000;
		color_arr[6908] = 8'b00001000;
		color_arr[6909] = 8'b00010010;
		color_arr[6910] = 8'b00010010;
		color_arr[6911] = 8'b00010010;
		color_arr[6912] = 8'b00010010;
		color_arr[6913] = 8'b00010010;
		color_arr[6914] = 8'b00000000;
		color_arr[6915] = 8'b00000000;
		color_arr[6916] = 8'b00010010;
		color_arr[6917] = 8'b00010010;
		color_arr[6918] = 8'b00010010;
		color_arr[6919] = 8'b00010010;
		color_arr[6920] = 8'b00000010;
		color_arr[6921] = 8'b00000010;
		color_arr[6922] = 8'b00000010;
		color_arr[6923] = 8'b00000010;
		color_arr[6924] = 8'b00000010;
		color_arr[6925] = 8'b00000010;
		color_arr[6926] = 8'b00000010;
		color_arr[6927] = 8'b00000010;
		color_arr[6928] = 8'b00000010;
		color_arr[6929] = 8'b00000010;
		color_arr[6930] = 8'b00000010;
		color_arr[6931] = 8'b00000010;
		color_arr[6932] = 8'b00000010;
		color_arr[6933] = 8'b00000010;
		color_arr[6934] = 8'b00000000;
		color_arr[6935] = 8'b00000000;
		color_arr[6936] = 8'b00000010;
		color_arr[6937] = 8'b00000010;
		color_arr[6938] = 8'b00000010;
		color_arr[6939] = 8'b00000010;
		color_arr[6940] = 8'b00000010;
		color_arr[6941] = 8'b00000010;
		color_arr[6942] = 8'b00000010;
		color_arr[6943] = 8'b00000010;
		color_arr[6944] = 8'b00000010;
		color_arr[6945] = 8'b00000010;
		color_arr[6946] = 8'b00000010;
		color_arr[6947] = 8'b00000010;
		color_arr[6948] = 8'b00000010;
		color_arr[6949] = 8'b00000010;
		color_arr[6950] = 8'b00100000;
		color_arr[6951] = 8'b00100000;
		color_arr[6952] = 8'b00100000;
		color_arr[6953] = 8'b00100000;
		color_arr[6954] = 8'b00100000;
		color_arr[6955] = 8'b00100000;
		color_arr[6956] = 8'b00100000;
		color_arr[6957] = 8'b00100000;
		color_arr[6958] = 8'b00100000;
		color_arr[6959] = 8'b00100000;
		color_arr[6960] = 8'b00100000;
		color_arr[6961] = 8'b00100000;
		color_arr[6962] = 8'b00100000;
		color_arr[6963] = 8'b00100000;
		color_arr[6964] = 8'b00100000;
		color_arr[6965] = 8'b00100000;
		color_arr[6966] = 8'b00100000;
		color_arr[6967] = 8'b00100000;
		color_arr[6968] = 8'b00100000;
		color_arr[6969] = 8'b00100000;
		color_arr[6970] = 8'b00100000;
		color_arr[6971] = 8'b00100000;
		color_arr[6972] = 8'b00100000;
		color_arr[6973] = 8'b00100000;
		color_arr[6974] = 8'b00100000;
		color_arr[6975] = 8'b00100000;
		color_arr[6976] = 8'b00100000;
		color_arr[6977] = 8'b00100000;
		color_arr[6978] = 8'b00100000;
		color_arr[6979] = 8'b00100000;
		color_arr[6980] = 8'b00100000;
		color_arr[6981] = 8'b00100000;
		color_arr[6982] = 8'b00100000;
		color_arr[6983] = 8'b00100000;
		color_arr[6984] = 8'b00100000;
		color_arr[6985] = 8'b00100000;
		color_arr[6986] = 8'b00100000;
		color_arr[6987] = 8'b00100000;
		color_arr[6988] = 8'b00100000;
		color_arr[6989] = 8'b00100000;
		color_arr[6990] = 8'b00100000;
		color_arr[6991] = 8'b00100000;
		color_arr[6992] = 8'b00001000;
		color_arr[6993] = 8'b00001000;
		color_arr[6994] = 8'b00001000;
		color_arr[6995] = 8'b00001000;
		color_arr[6996] = 8'b00001000;
		color_arr[6997] = 8'b00001000;
		color_arr[6998] = 8'b00001000;
		color_arr[6999] = 8'b00001000;
		color_arr[7000] = 8'b00001000;
		color_arr[7001] = 8'b00001000;
		color_arr[7002] = 8'b00001000;
		color_arr[7003] = 8'b00001000;
		color_arr[7004] = 8'b00001000;
		color_arr[7005] = 8'b00001000;
		color_arr[7006] = 8'b00001000;
		color_arr[7007] = 8'b00001000;
		color_arr[7008] = 8'b00000000;
		color_arr[7009] = 8'b00000000;
		color_arr[7010] = 8'b00001000;
		color_arr[7011] = 8'b00001000;
		color_arr[7012] = 8'b00001000;
		color_arr[7013] = 8'b00001000;
		color_arr[7014] = 8'b00001000;
		color_arr[7015] = 8'b00001000;
		color_arr[7016] = 8'b00001000;
		color_arr[7017] = 8'b00001000;
		color_arr[7018] = 8'b00001000;
		color_arr[7019] = 8'b00000000;
		color_arr[7020] = 8'b00000000;
		color_arr[7021] = 8'b00000000;
		color_arr[7022] = 8'b00001000;
		color_arr[7023] = 8'b00001000;
		color_arr[7024] = 8'b00001000;
		color_arr[7025] = 8'b00001000;
		color_arr[7026] = 8'b00001000;
		color_arr[7027] = 8'b00001000;
		color_arr[7028] = 8'b00000000;
		color_arr[7029] = 8'b00000000;
		color_arr[7030] = 8'b00001000;
		color_arr[7031] = 8'b00001000;
		color_arr[7032] = 8'b00001000;
		color_arr[7033] = 8'b00001000;
		color_arr[7034] = 8'b00001000;
		color_arr[7035] = 8'b00001000;
		color_arr[7036] = 8'b00001000;
		color_arr[7037] = 8'b00010010;
		color_arr[7038] = 8'b00010010;
		color_arr[7039] = 8'b00010010;
		color_arr[7040] = 8'b00010010;
		color_arr[7041] = 8'b00010010;
		color_arr[7042] = 8'b00000000;
		color_arr[7043] = 8'b00000000;
		color_arr[7044] = 8'b00010010;
		color_arr[7045] = 8'b00010010;
		color_arr[7046] = 8'b00010010;
		color_arr[7047] = 8'b00010010;
		color_arr[7048] = 8'b00010010;
		color_arr[7049] = 8'b00010010;
		color_arr[7050] = 8'b00010010;
		color_arr[7051] = 8'b00010010;
		color_arr[7052] = 8'b00010010;
		color_arr[7053] = 8'b00010010;
		color_arr[7054] = 8'b00010010;
		color_arr[7055] = 8'b00010010;
		color_arr[7056] = 8'b00010010;
		color_arr[7057] = 8'b00010010;
		color_arr[7058] = 8'b00100000;
		color_arr[7059] = 8'b00100000;
		color_arr[7060] = 8'b00100000;
		color_arr[7061] = 8'b00100000;
		color_arr[7062] = 8'b00000000;
		color_arr[7063] = 8'b00000000;
		color_arr[7064] = 8'b00100000;
		color_arr[7065] = 8'b00100000;
		color_arr[7066] = 8'b00100000;
		color_arr[7067] = 8'b00100000;
		color_arr[7068] = 8'b00100000;
		color_arr[7069] = 8'b00100000;
		color_arr[7070] = 8'b00100000;
		color_arr[7071] = 8'b00100000;
		color_arr[7072] = 8'b00100000;
		color_arr[7073] = 8'b00100000;
		color_arr[7074] = 8'b00100000;
		color_arr[7075] = 8'b00100000;
		color_arr[7076] = 8'b00100000;
		color_arr[7077] = 8'b00100000;
		color_arr[7078] = 8'b00100000;
		color_arr[7079] = 8'b00100000;
		color_arr[7080] = 8'b00100000;
		color_arr[7081] = 8'b00100000;
		color_arr[7082] = 8'b00100000;
		color_arr[7083] = 8'b00100000;
		color_arr[7084] = 8'b00100000;
		color_arr[7085] = 8'b00100000;
		color_arr[7086] = 8'b00100000;
		color_arr[7087] = 8'b00100000;
		color_arr[7088] = 8'b00100000;
		color_arr[7089] = 8'b00100000;
		color_arr[7090] = 8'b00100000;
		color_arr[7091] = 8'b00100000;
		color_arr[7092] = 8'b00100000;
		color_arr[7093] = 8'b00100000;
		color_arr[7094] = 8'b00100000;
		color_arr[7095] = 8'b00100000;
		color_arr[7096] = 8'b00100000;
		color_arr[7097] = 8'b00100000;
		color_arr[7098] = 8'b00100000;
		color_arr[7099] = 8'b00100000;
		color_arr[7100] = 8'b00100000;
		color_arr[7101] = 8'b00100000;
		color_arr[7102] = 8'b00100000;
		color_arr[7103] = 8'b00100000;
		color_arr[7104] = 8'b00100000;
		color_arr[7105] = 8'b00100000;
		color_arr[7106] = 8'b00100000;
		color_arr[7107] = 8'b00100000;
		color_arr[7108] = 8'b00100000;
		color_arr[7109] = 8'b00100000;
		color_arr[7110] = 8'b00100000;
		color_arr[7111] = 8'b00100000;
		color_arr[7112] = 8'b00100000;
		color_arr[7113] = 8'b00100000;
		color_arr[7114] = 8'b00100000;
		color_arr[7115] = 8'b00100000;
		color_arr[7116] = 8'b00100000;
		color_arr[7117] = 8'b00100000;
		color_arr[7118] = 8'b00100000;
		color_arr[7119] = 8'b00100000;
		color_arr[7120] = 8'b00001000;
		color_arr[7121] = 8'b00001000;
		color_arr[7122] = 8'b00001000;
		color_arr[7123] = 8'b00001000;
		color_arr[7124] = 8'b00001000;
		color_arr[7125] = 8'b00001000;
		color_arr[7126] = 8'b00001000;
		color_arr[7127] = 8'b00001000;
		color_arr[7128] = 8'b00001000;
		color_arr[7129] = 8'b00001000;
		color_arr[7130] = 8'b00001000;
		color_arr[7131] = 8'b00001000;
		color_arr[7132] = 8'b00001000;
		color_arr[7133] = 8'b00001000;
		color_arr[7134] = 8'b00001000;
		color_arr[7135] = 8'b00001000;
		color_arr[7136] = 8'b00000000;
		color_arr[7137] = 8'b00000000;
		color_arr[7138] = 8'b00001000;
		color_arr[7139] = 8'b00001000;
		color_arr[7140] = 8'b00001000;
		color_arr[7141] = 8'b00001000;
		color_arr[7142] = 8'b00001000;
		color_arr[7143] = 8'b00001000;
		color_arr[7144] = 8'b00001000;
		color_arr[7145] = 8'b00001000;
		color_arr[7146] = 8'b00001000;
		color_arr[7147] = 8'b00001000;
		color_arr[7148] = 8'b00000000;
		color_arr[7149] = 8'b00000000;
		color_arr[7150] = 8'b00000000;
		color_arr[7151] = 8'b00001000;
		color_arr[7152] = 8'b00001000;
		color_arr[7153] = 8'b00001000;
		color_arr[7154] = 8'b00001000;
		color_arr[7155] = 8'b00001000;
		color_arr[7156] = 8'b00000000;
		color_arr[7157] = 8'b00000000;
		color_arr[7158] = 8'b00001000;
		color_arr[7159] = 8'b00001000;
		color_arr[7160] = 8'b00001000;
		color_arr[7161] = 8'b00001000;
		color_arr[7162] = 8'b00001000;
		color_arr[7163] = 8'b00001000;
		color_arr[7164] = 8'b00001000;
		color_arr[7165] = 8'b00010010;
		color_arr[7166] = 8'b00010010;
		color_arr[7167] = 8'b00010010;
		color_arr[7168] = 8'b00010010;
		color_arr[7169] = 8'b00010010;
		color_arr[7170] = 8'b00000000;
		color_arr[7171] = 8'b00000000;
		color_arr[7172] = 8'b00010010;
		color_arr[7173] = 8'b00010010;
		color_arr[7174] = 8'b00010010;
		color_arr[7175] = 8'b00010010;
		color_arr[7176] = 8'b00010010;
		color_arr[7177] = 8'b00010010;
		color_arr[7178] = 8'b00010010;
		color_arr[7179] = 8'b00010010;
		color_arr[7180] = 8'b00010010;
		color_arr[7181] = 8'b00010010;
		color_arr[7182] = 8'b00010010;
		color_arr[7183] = 8'b00010010;
		color_arr[7184] = 8'b00010010;
		color_arr[7185] = 8'b00010010;
		color_arr[7186] = 8'b00100000;
		color_arr[7187] = 8'b00100000;
		color_arr[7188] = 8'b00100000;
		color_arr[7189] = 8'b00000000;
		color_arr[7190] = 8'b00000000;
		color_arr[7191] = 8'b00000000;
		color_arr[7192] = 8'b00100000;
		color_arr[7193] = 8'b00100000;
		color_arr[7194] = 8'b00100000;
		color_arr[7195] = 8'b00100000;
		color_arr[7196] = 8'b00100000;
		color_arr[7197] = 8'b00100000;
		color_arr[7198] = 8'b00100000;
		color_arr[7199] = 8'b00100000;
		color_arr[7200] = 8'b00100000;
		color_arr[7201] = 8'b00100000;
		color_arr[7202] = 8'b00100000;
		color_arr[7203] = 8'b00100000;
		color_arr[7204] = 8'b00100000;
		color_arr[7205] = 8'b00100000;
		color_arr[7206] = 8'b00100000;
		color_arr[7207] = 8'b00100000;
		color_arr[7208] = 8'b00100000;
		color_arr[7209] = 8'b00100000;
		color_arr[7210] = 8'b00100000;
		color_arr[7211] = 8'b00100000;
		color_arr[7212] = 8'b00100000;
		color_arr[7213] = 8'b00100000;
		color_arr[7214] = 8'b00100000;
		color_arr[7215] = 8'b00100000;
		color_arr[7216] = 8'b00100000;
		color_arr[7217] = 8'b00100000;
		color_arr[7218] = 8'b00100000;
		color_arr[7219] = 8'b00100000;
		color_arr[7220] = 8'b00100000;
		color_arr[7221] = 8'b00100000;
		color_arr[7222] = 8'b00100000;
		color_arr[7223] = 8'b00100000;
		color_arr[7224] = 8'b00100000;
		color_arr[7225] = 8'b00100000;
		color_arr[7226] = 8'b00100000;
		color_arr[7227] = 8'b00100000;
		color_arr[7228] = 8'b00100000;
		color_arr[7229] = 8'b00100000;
		color_arr[7230] = 8'b00100000;
		color_arr[7231] = 8'b00100000;
		color_arr[7232] = 8'b00100000;
		color_arr[7233] = 8'b00100000;
		color_arr[7234] = 8'b00100000;
		color_arr[7235] = 8'b00100000;
		color_arr[7236] = 8'b00100000;
		color_arr[7237] = 8'b00100000;
		color_arr[7238] = 8'b00100000;
		color_arr[7239] = 8'b00100000;
		color_arr[7240] = 8'b00100000;
		color_arr[7241] = 8'b00100000;
		color_arr[7242] = 8'b00100000;
		color_arr[7243] = 8'b00100000;
		color_arr[7244] = 8'b00100000;
		color_arr[7245] = 8'b00100000;
		color_arr[7246] = 8'b00100000;
		color_arr[7247] = 8'b00100000;
		color_arr[7248] = 8'b00001000;
		color_arr[7249] = 8'b00001000;
		color_arr[7250] = 8'b00001000;
		color_arr[7251] = 8'b00001000;
		color_arr[7252] = 8'b00001000;
		color_arr[7253] = 8'b00001000;
		color_arr[7254] = 8'b00001000;
		color_arr[7255] = 8'b00001000;
		color_arr[7256] = 8'b00001000;
		color_arr[7257] = 8'b00001000;
		color_arr[7258] = 8'b00001000;
		color_arr[7259] = 8'b00001000;
		color_arr[7260] = 8'b00001000;
		color_arr[7261] = 8'b00001000;
		color_arr[7262] = 8'b00001000;
		color_arr[7263] = 8'b00000000;
		color_arr[7264] = 8'b00000000;
		color_arr[7265] = 8'b00000000;
		color_arr[7266] = 8'b00001000;
		color_arr[7267] = 8'b00001000;
		color_arr[7268] = 8'b00001000;
		color_arr[7269] = 8'b00001000;
		color_arr[7270] = 8'b00001000;
		color_arr[7271] = 8'b00001000;
		color_arr[7272] = 8'b00001000;
		color_arr[7273] = 8'b00001000;
		color_arr[7274] = 8'b00001000;
		color_arr[7275] = 8'b00001000;
		color_arr[7276] = 8'b00001000;
		color_arr[7277] = 8'b00000000;
		color_arr[7278] = 8'b00000000;
		color_arr[7279] = 8'b00001000;
		color_arr[7280] = 8'b00001000;
		color_arr[7281] = 8'b00001000;
		color_arr[7282] = 8'b00001000;
		color_arr[7283] = 8'b00001000;
		color_arr[7284] = 8'b00000000;
		color_arr[7285] = 8'b00000000;
		color_arr[7286] = 8'b00001000;
		color_arr[7287] = 8'b00001000;
		color_arr[7288] = 8'b00001000;
		color_arr[7289] = 8'b00001000;
		color_arr[7290] = 8'b00001000;
		color_arr[7291] = 8'b00001000;
		color_arr[7292] = 8'b00001000;
		color_arr[7293] = 8'b00010010;
		color_arr[7294] = 8'b00010010;
		color_arr[7295] = 8'b00010010;
		color_arr[7296] = 8'b00010010;
		color_arr[7297] = 8'b00010010;
		color_arr[7298] = 8'b00000000;
		color_arr[7299] = 8'b00000000;
		color_arr[7300] = 8'b00010010;
		color_arr[7301] = 8'b00010010;
		color_arr[7302] = 8'b00010010;
		color_arr[7303] = 8'b00010010;
		color_arr[7304] = 8'b00010010;
		color_arr[7305] = 8'b00010010;
		color_arr[7306] = 8'b00010010;
		color_arr[7307] = 8'b00010010;
		color_arr[7308] = 8'b00010010;
		color_arr[7309] = 8'b00010010;
		color_arr[7310] = 8'b00010010;
		color_arr[7311] = 8'b00010010;
		color_arr[7312] = 8'b00010010;
		color_arr[7313] = 8'b00010010;
		color_arr[7314] = 8'b00100000;
		color_arr[7315] = 8'b00100000;
		color_arr[7316] = 8'b00100000;
		color_arr[7317] = 8'b00000000;
		color_arr[7318] = 8'b00000000;
		color_arr[7319] = 8'b00100000;
		color_arr[7320] = 8'b00100000;
		color_arr[7321] = 8'b00100000;
		color_arr[7322] = 8'b00100000;
		color_arr[7323] = 8'b00100000;
		color_arr[7324] = 8'b00100000;
		color_arr[7325] = 8'b00100000;
		color_arr[7326] = 8'b00100000;
		color_arr[7327] = 8'b00100000;
		color_arr[7328] = 8'b00100000;
		color_arr[7329] = 8'b00100000;
		color_arr[7330] = 8'b00100000;
		color_arr[7331] = 8'b00100000;
		color_arr[7332] = 8'b00100000;
		color_arr[7333] = 8'b00100000;
		color_arr[7334] = 8'b00100000;
		color_arr[7335] = 8'b00100000;
		color_arr[7336] = 8'b00100000;
		color_arr[7337] = 8'b00100000;
		color_arr[7338] = 8'b00100000;
		color_arr[7339] = 8'b00100000;
		color_arr[7340] = 8'b00100000;
		color_arr[7341] = 8'b00100000;
		color_arr[7342] = 8'b00100000;
		color_arr[7343] = 8'b00100000;
		color_arr[7344] = 8'b00100000;
		color_arr[7345] = 8'b00100000;
		color_arr[7346] = 8'b00100000;
		color_arr[7347] = 8'b00100000;
		color_arr[7348] = 8'b00100000;
		color_arr[7349] = 8'b00100000;
		color_arr[7350] = 8'b00100000;
		color_arr[7351] = 8'b00100000;
		color_arr[7352] = 8'b00100000;
		color_arr[7353] = 8'b00100000;
		color_arr[7354] = 8'b00100000;
		color_arr[7355] = 8'b00100000;
		color_arr[7356] = 8'b00100000;
		color_arr[7357] = 8'b00100000;
		color_arr[7358] = 8'b00100000;
		color_arr[7359] = 8'b00100000;
		color_arr[7360] = 8'b00100000;
		color_arr[7361] = 8'b00100000;
		color_arr[7362] = 8'b00100000;
		color_arr[7363] = 8'b00100000;
		color_arr[7364] = 8'b00100000;
		color_arr[7365] = 8'b00100000;
		color_arr[7366] = 8'b00100000;
		color_arr[7367] = 8'b00100000;
		color_arr[7368] = 8'b00100000;
		color_arr[7369] = 8'b00100000;
		color_arr[7370] = 8'b00100000;
		color_arr[7371] = 8'b00100000;
		color_arr[7372] = 8'b00100000;
		color_arr[7373] = 8'b00100000;
		color_arr[7374] = 8'b00100000;
		color_arr[7375] = 8'b00100000;
		color_arr[7376] = 8'b00001000;
		color_arr[7377] = 8'b00001000;
		color_arr[7378] = 8'b00001000;
		color_arr[7379] = 8'b00001000;
		color_arr[7380] = 8'b00001000;
		color_arr[7381] = 8'b00001000;
		color_arr[7382] = 8'b00001000;
		color_arr[7383] = 8'b00001000;
		color_arr[7384] = 8'b00001000;
		color_arr[7385] = 8'b00001000;
		color_arr[7386] = 8'b00001000;
		color_arr[7387] = 8'b00001000;
		color_arr[7388] = 8'b00001000;
		color_arr[7389] = 8'b00001000;
		color_arr[7390] = 8'b00001000;
		color_arr[7391] = 8'b00000000;
		color_arr[7392] = 8'b00000000;
		color_arr[7393] = 8'b00001000;
		color_arr[7394] = 8'b00001000;
		color_arr[7395] = 8'b00001000;
		color_arr[7396] = 8'b00001000;
		color_arr[7397] = 8'b00001000;
		color_arr[7398] = 8'b00001000;
		color_arr[7399] = 8'b00001000;
		color_arr[7400] = 8'b00001000;
		color_arr[7401] = 8'b00001000;
		color_arr[7402] = 8'b00001000;
		color_arr[7403] = 8'b00001000;
		color_arr[7404] = 8'b00001000;
		color_arr[7405] = 8'b00000000;
		color_arr[7406] = 8'b00000000;
		color_arr[7407] = 8'b00000000;
		color_arr[7408] = 8'b00001000;
		color_arr[7409] = 8'b00001000;
		color_arr[7410] = 8'b00001000;
		color_arr[7411] = 8'b00001000;
		color_arr[7412] = 8'b00000000;
		color_arr[7413] = 8'b00000000;
		color_arr[7414] = 8'b00001000;
		color_arr[7415] = 8'b00001000;
		color_arr[7416] = 8'b00001000;
		color_arr[7417] = 8'b00001000;
		color_arr[7418] = 8'b00001000;
		color_arr[7419] = 8'b00001000;
		color_arr[7420] = 8'b00001000;
		color_arr[7421] = 8'b00010010;
		color_arr[7422] = 8'b00010010;
		color_arr[7423] = 8'b00010010;
		color_arr[7424] = 8'b00010010;
		color_arr[7425] = 8'b00010010;
		color_arr[7426] = 8'b00000000;
		color_arr[7427] = 8'b00000000;
		color_arr[7428] = 8'b00010010;
		color_arr[7429] = 8'b00010010;
		color_arr[7430] = 8'b00010010;
		color_arr[7431] = 8'b00010010;
		color_arr[7432] = 8'b00010010;
		color_arr[7433] = 8'b00010010;
		color_arr[7434] = 8'b00010010;
		color_arr[7435] = 8'b00010010;
		color_arr[7436] = 8'b00010010;
		color_arr[7437] = 8'b00010010;
		color_arr[7438] = 8'b00010010;
		color_arr[7439] = 8'b00010010;
		color_arr[7440] = 8'b00010010;
		color_arr[7441] = 8'b00010010;
		color_arr[7442] = 8'b00100000;
		color_arr[7443] = 8'b00100000;
		color_arr[7444] = 8'b00100000;
		color_arr[7445] = 8'b00000000;
		color_arr[7446] = 8'b00000000;
		color_arr[7447] = 8'b00100000;
		color_arr[7448] = 8'b00100000;
		color_arr[7449] = 8'b00100000;
		color_arr[7450] = 8'b00100000;
		color_arr[7451] = 8'b00100000;
		color_arr[7452] = 8'b00100000;
		color_arr[7453] = 8'b00100000;
		color_arr[7454] = 8'b00100000;
		color_arr[7455] = 8'b00100000;
		color_arr[7456] = 8'b00100000;
		color_arr[7457] = 8'b00100000;
		color_arr[7458] = 8'b00100000;
		color_arr[7459] = 8'b00100000;
		color_arr[7460] = 8'b00100000;
		color_arr[7461] = 8'b00100000;
		color_arr[7462] = 8'b00100000;
		color_arr[7463] = 8'b00100000;
		color_arr[7464] = 8'b00100000;
		color_arr[7465] = 8'b00100000;
		color_arr[7466] = 8'b00100000;
		color_arr[7467] = 8'b00100000;
		color_arr[7468] = 8'b00100000;
		color_arr[7469] = 8'b00100000;
		color_arr[7470] = 8'b00100000;
		color_arr[7471] = 8'b00100000;
		color_arr[7472] = 8'b00100000;
		color_arr[7473] = 8'b00100000;
		color_arr[7474] = 8'b00100000;
		color_arr[7475] = 8'b00100000;
		color_arr[7476] = 8'b00100000;
		color_arr[7477] = 8'b00100000;
		color_arr[7478] = 8'b00100000;
		color_arr[7479] = 8'b00100000;
		color_arr[7480] = 8'b00100000;
		color_arr[7481] = 8'b00100000;
		color_arr[7482] = 8'b00100000;
		color_arr[7483] = 8'b00100000;
		color_arr[7484] = 8'b00100000;
		color_arr[7485] = 8'b00100000;
		color_arr[7486] = 8'b00100000;
		color_arr[7487] = 8'b00100000;
		color_arr[7488] = 8'b00100000;
		color_arr[7489] = 8'b00100000;
		color_arr[7490] = 8'b00100000;
		color_arr[7491] = 8'b00100000;
		color_arr[7492] = 8'b00100000;
		color_arr[7493] = 8'b00100000;
		color_arr[7494] = 8'b00100000;
		color_arr[7495] = 8'b00100000;
		color_arr[7496] = 8'b00100000;
		color_arr[7497] = 8'b00100000;
		color_arr[7498] = 8'b00100000;
		color_arr[7499] = 8'b00100000;
		color_arr[7500] = 8'b00100000;
		color_arr[7501] = 8'b00100000;
		color_arr[7502] = 8'b00100000;
		color_arr[7503] = 8'b00100000;
		color_arr[7504] = 8'b00001000;
		color_arr[7505] = 8'b00001000;
		color_arr[7506] = 8'b00001000;
		color_arr[7507] = 8'b00001000;
		color_arr[7508] = 8'b00001000;
		color_arr[7509] = 8'b00001000;
		color_arr[7510] = 8'b00001000;
		color_arr[7511] = 8'b00001000;
		color_arr[7512] = 8'b00001000;
		color_arr[7513] = 8'b00001000;
		color_arr[7514] = 8'b00001000;
		color_arr[7515] = 8'b00001000;
		color_arr[7516] = 8'b00001000;
		color_arr[7517] = 8'b00001000;
		color_arr[7518] = 8'b00000000;
		color_arr[7519] = 8'b00000000;
		color_arr[7520] = 8'b00000000;
		color_arr[7521] = 8'b00001000;
		color_arr[7522] = 8'b00001000;
		color_arr[7523] = 8'b00001000;
		color_arr[7524] = 8'b00001000;
		color_arr[7525] = 8'b00001000;
		color_arr[7526] = 8'b00001000;
		color_arr[7527] = 8'b00001000;
		color_arr[7528] = 8'b00001000;
		color_arr[7529] = 8'b00001000;
		color_arr[7530] = 8'b00001000;
		color_arr[7531] = 8'b00001000;
		color_arr[7532] = 8'b00001000;
		color_arr[7533] = 8'b00001000;
		color_arr[7534] = 8'b00000000;
		color_arr[7535] = 8'b00000000;
		color_arr[7536] = 8'b00001000;
		color_arr[7537] = 8'b00001000;
		color_arr[7538] = 8'b00001000;
		color_arr[7539] = 8'b00001000;
		color_arr[7540] = 8'b00000000;
		color_arr[7541] = 8'b00000000;
		color_arr[7542] = 8'b00001000;
		color_arr[7543] = 8'b00001000;
		color_arr[7544] = 8'b00001000;
		color_arr[7545] = 8'b00001000;
		color_arr[7546] = 8'b00001000;
		color_arr[7547] = 8'b00001000;
		color_arr[7548] = 8'b00001000;
		color_arr[7549] = 8'b00010010;
		color_arr[7550] = 8'b00010010;
		color_arr[7551] = 8'b00010010;
		color_arr[7552] = 8'b00010010;
		color_arr[7553] = 8'b00010010;
		color_arr[7554] = 8'b00000000;
		color_arr[7555] = 8'b00000000;
		color_arr[7556] = 8'b00010010;
		color_arr[7557] = 8'b00010010;
		color_arr[7558] = 8'b00010010;
		color_arr[7559] = 8'b00010010;
		color_arr[7560] = 8'b00010010;
		color_arr[7561] = 8'b00010010;
		color_arr[7562] = 8'b00010010;
		color_arr[7563] = 8'b00010010;
		color_arr[7564] = 8'b00010010;
		color_arr[7565] = 8'b00010010;
		color_arr[7566] = 8'b00010010;
		color_arr[7567] = 8'b00010010;
		color_arr[7568] = 8'b00010010;
		color_arr[7569] = 8'b00010010;
		color_arr[7570] = 8'b00100000;
		color_arr[7571] = 8'b00100000;
		color_arr[7572] = 8'b00100000;
		color_arr[7573] = 8'b00000000;
		color_arr[7574] = 8'b00000000;
		color_arr[7575] = 8'b00100000;
		color_arr[7576] = 8'b00100000;
		color_arr[7577] = 8'b00100000;
		color_arr[7578] = 8'b00100000;
		color_arr[7579] = 8'b00100000;
		color_arr[7580] = 8'b00100000;
		color_arr[7581] = 8'b00100000;
		color_arr[7582] = 8'b00100000;
		color_arr[7583] = 8'b00100000;
		color_arr[7584] = 8'b00100000;
		color_arr[7585] = 8'b00100000;
		color_arr[7586] = 8'b00100000;
		color_arr[7587] = 8'b00100000;
		color_arr[7588] = 8'b00100000;
		color_arr[7589] = 8'b00100000;
		color_arr[7590] = 8'b00100000;
		color_arr[7591] = 8'b00100000;
		color_arr[7592] = 8'b00100000;
		color_arr[7593] = 8'b00100000;
		color_arr[7594] = 8'b00100000;
		color_arr[7595] = 8'b00100000;
		color_arr[7596] = 8'b00100000;
		color_arr[7597] = 8'b00100000;
		color_arr[7598] = 8'b00100000;
		color_arr[7599] = 8'b00100000;
		color_arr[7600] = 8'b00100000;
		color_arr[7601] = 8'b00100000;
		color_arr[7602] = 8'b00100000;
		color_arr[7603] = 8'b00100000;
		color_arr[7604] = 8'b00100000;
		color_arr[7605] = 8'b00100000;
		color_arr[7606] = 8'b00100000;
		color_arr[7607] = 8'b00100000;
		color_arr[7608] = 8'b00100000;
		color_arr[7609] = 8'b00100000;
		color_arr[7610] = 8'b00100000;
		color_arr[7611] = 8'b00100000;
		color_arr[7612] = 8'b00100000;
		color_arr[7613] = 8'b00100000;
		color_arr[7614] = 8'b00100000;
		color_arr[7615] = 8'b00100000;
		color_arr[7616] = 8'b00100000;
		color_arr[7617] = 8'b00100000;
		color_arr[7618] = 8'b00100000;
		color_arr[7619] = 8'b00100000;
		color_arr[7620] = 8'b00100000;
		color_arr[7621] = 8'b00100000;
		color_arr[7622] = 8'b00100000;
		color_arr[7623] = 8'b00100000;
		color_arr[7624] = 8'b00100000;
		color_arr[7625] = 8'b00100000;
		color_arr[7626] = 8'b00100000;
		color_arr[7627] = 8'b00100000;
		color_arr[7628] = 8'b00100000;
		color_arr[7629] = 8'b00100000;
		color_arr[7630] = 8'b00100000;
		color_arr[7631] = 8'b00100000;
		color_arr[7632] = 8'b00001000;
		color_arr[7633] = 8'b00001000;
		color_arr[7634] = 8'b00001000;
		color_arr[7635] = 8'b00001000;
		color_arr[7636] = 8'b00001000;
		color_arr[7637] = 8'b00001000;
		color_arr[7638] = 8'b00001000;
		color_arr[7639] = 8'b00001000;
		color_arr[7640] = 8'b00001000;
		color_arr[7641] = 8'b00001000;
		color_arr[7642] = 8'b00001000;
		color_arr[7643] = 8'b00001000;
		color_arr[7644] = 8'b00001000;
		color_arr[7645] = 8'b00001000;
		color_arr[7646] = 8'b00000000;
		color_arr[7647] = 8'b00000000;
		color_arr[7648] = 8'b00001000;
		color_arr[7649] = 8'b00001000;
		color_arr[7650] = 8'b00001000;
		color_arr[7651] = 8'b00001000;
		color_arr[7652] = 8'b00001000;
		color_arr[7653] = 8'b00001000;
		color_arr[7654] = 8'b00001000;
		color_arr[7655] = 8'b00001000;
		color_arr[7656] = 8'b00001000;
		color_arr[7657] = 8'b00001000;
		color_arr[7658] = 8'b00001000;
		color_arr[7659] = 8'b00001000;
		color_arr[7660] = 8'b00001000;
		color_arr[7661] = 8'b00001000;
		color_arr[7662] = 8'b00000000;
		color_arr[7663] = 8'b00000000;
		color_arr[7664] = 8'b00000000;
		color_arr[7665] = 8'b00001000;
		color_arr[7666] = 8'b00001000;
		color_arr[7667] = 8'b00001000;
		color_arr[7668] = 8'b00000000;
		color_arr[7669] = 8'b00000000;
		color_arr[7670] = 8'b00001000;
		color_arr[7671] = 8'b00001000;
		color_arr[7672] = 8'b00001000;
		color_arr[7673] = 8'b00001000;
		color_arr[7674] = 8'b00001000;
		color_arr[7675] = 8'b00001000;
		color_arr[7676] = 8'b00001000;
		color_arr[7677] = 8'b00010010;
		color_arr[7678] = 8'b00010010;
		color_arr[7679] = 8'b00010010;
		color_arr[7680] = 8'b00010010;
		color_arr[7681] = 8'b00010010;
		color_arr[7682] = 8'b00000000;
		color_arr[7683] = 8'b00000000;
		color_arr[7684] = 8'b00010010;
		color_arr[7685] = 8'b00010010;
		color_arr[7686] = 8'b00010010;
		color_arr[7687] = 8'b00010010;
		color_arr[7688] = 8'b00010010;
		color_arr[7689] = 8'b00010010;
		color_arr[7690] = 8'b00010010;
		color_arr[7691] = 8'b00010010;
		color_arr[7692] = 8'b00010010;
		color_arr[7693] = 8'b00010010;
		color_arr[7694] = 8'b00010010;
		color_arr[7695] = 8'b00010010;
		color_arr[7696] = 8'b00010010;
		color_arr[7697] = 8'b00010010;
		color_arr[7698] = 8'b00100000;
		color_arr[7699] = 8'b00100000;
		color_arr[7700] = 8'b00100000;
		color_arr[7701] = 8'b00000000;
		color_arr[7702] = 8'b00000000;
		color_arr[7703] = 8'b00100000;
		color_arr[7704] = 8'b00100000;
		color_arr[7705] = 8'b00100000;
		color_arr[7706] = 8'b00100000;
		color_arr[7707] = 8'b00100000;
		color_arr[7708] = 8'b00100000;
		color_arr[7709] = 8'b00100000;
		color_arr[7710] = 8'b00100000;
		color_arr[7711] = 8'b00100000;
		color_arr[7712] = 8'b00100000;
		color_arr[7713] = 8'b00100000;
		color_arr[7714] = 8'b00100000;
		color_arr[7715] = 8'b00100000;
		color_arr[7716] = 8'b00100000;
		color_arr[7717] = 8'b00100000;
		color_arr[7718] = 8'b00100000;
		color_arr[7719] = 8'b00100000;
		color_arr[7720] = 8'b00100000;
		color_arr[7721] = 8'b00100000;
		color_arr[7722] = 8'b00100000;
		color_arr[7723] = 8'b00100000;
		color_arr[7724] = 8'b00100000;
		color_arr[7725] = 8'b00100000;
		color_arr[7726] = 8'b00100000;
		color_arr[7727] = 8'b00100000;
		color_arr[7728] = 8'b00100000;
		color_arr[7729] = 8'b00100000;
		color_arr[7730] = 8'b00100000;
		color_arr[7731] = 8'b00100000;
		color_arr[7732] = 8'b00100000;
		color_arr[7733] = 8'b00100000;
		color_arr[7734] = 8'b00100000;
		color_arr[7735] = 8'b00100000;
		color_arr[7736] = 8'b00100000;
		color_arr[7737] = 8'b00100000;
		color_arr[7738] = 8'b00100000;
		color_arr[7739] = 8'b00100000;
		color_arr[7740] = 8'b00100000;
		color_arr[7741] = 8'b00100000;
		color_arr[7742] = 8'b00100000;
		color_arr[7743] = 8'b00100000;
		color_arr[7744] = 8'b00100000;
		color_arr[7745] = 8'b00100000;
		color_arr[7746] = 8'b00100000;
		color_arr[7747] = 8'b00100000;
		color_arr[7748] = 8'b00100000;
		color_arr[7749] = 8'b00100000;
		color_arr[7750] = 8'b00100000;
		color_arr[7751] = 8'b00100000;
		color_arr[7752] = 8'b00100000;
		color_arr[7753] = 8'b00100000;
		color_arr[7754] = 8'b00100000;
		color_arr[7755] = 8'b00100000;
		color_arr[7756] = 8'b00100000;
		color_arr[7757] = 8'b00100000;
		color_arr[7758] = 8'b00100000;
		color_arr[7759] = 8'b00100000;
		color_arr[7760] = 8'b00001000;
		color_arr[7761] = 8'b00001000;
		color_arr[7762] = 8'b00001000;
		color_arr[7763] = 8'b00001000;
		color_arr[7764] = 8'b00001000;
		color_arr[7765] = 8'b00001000;
		color_arr[7766] = 8'b00001000;
		color_arr[7767] = 8'b00001000;
		color_arr[7768] = 8'b00001000;
		color_arr[7769] = 8'b00001000;
		color_arr[7770] = 8'b00001000;
		color_arr[7771] = 8'b00001000;
		color_arr[7772] = 8'b00001000;
		color_arr[7773] = 8'b00000000;
		color_arr[7774] = 8'b00000000;
		color_arr[7775] = 8'b00000000;
		color_arr[7776] = 8'b00001000;
		color_arr[7777] = 8'b00001000;
		color_arr[7778] = 8'b00001000;
		color_arr[7779] = 8'b00001000;
		color_arr[7780] = 8'b00001000;
		color_arr[7781] = 8'b00001000;
		color_arr[7782] = 8'b00001000;
		color_arr[7783] = 8'b00001000;
		color_arr[7784] = 8'b00001000;
		color_arr[7785] = 8'b00001000;
		color_arr[7786] = 8'b00001000;
		color_arr[7787] = 8'b00001000;
		color_arr[7788] = 8'b00001000;
		color_arr[7789] = 8'b00001000;
		color_arr[7790] = 8'b00001000;
		color_arr[7791] = 8'b00000000;
		color_arr[7792] = 8'b00000000;
		color_arr[7793] = 8'b00001000;
		color_arr[7794] = 8'b00001000;
		color_arr[7795] = 8'b00001000;
		color_arr[7796] = 8'b00000000;
		color_arr[7797] = 8'b00000000;
		color_arr[7798] = 8'b00000000;
		color_arr[7799] = 8'b00001000;
		color_arr[7800] = 8'b00001000;
		color_arr[7801] = 8'b00001000;
		color_arr[7802] = 8'b00001000;
		color_arr[7803] = 8'b00001000;
		color_arr[7804] = 8'b00001000;
		color_arr[7805] = 8'b00010010;
		color_arr[7806] = 8'b00010010;
		color_arr[7807] = 8'b00010010;
		color_arr[7808] = 8'b00010010;
		color_arr[7809] = 8'b00010010;
		color_arr[7810] = 8'b00000000;
		color_arr[7811] = 8'b00000000;
		color_arr[7812] = 8'b00010010;
		color_arr[7813] = 8'b00010010;
		color_arr[7814] = 8'b00010010;
		color_arr[7815] = 8'b00010010;
		color_arr[7816] = 8'b00010010;
		color_arr[7817] = 8'b00010010;
		color_arr[7818] = 8'b00010010;
		color_arr[7819] = 8'b00010010;
		color_arr[7820] = 8'b00010010;
		color_arr[7821] = 8'b00010010;
		color_arr[7822] = 8'b00010010;
		color_arr[7823] = 8'b00010010;
		color_arr[7824] = 8'b00010010;
		color_arr[7825] = 8'b00010010;
		color_arr[7826] = 8'b00100000;
		color_arr[7827] = 8'b00100000;
		color_arr[7828] = 8'b00100000;
		color_arr[7829] = 8'b00000000;
		color_arr[7830] = 8'b00000000;
		color_arr[7831] = 8'b00100000;
		color_arr[7832] = 8'b00100000;
		color_arr[7833] = 8'b00100000;
		color_arr[7834] = 8'b00100000;
		color_arr[7835] = 8'b00100000;
		color_arr[7836] = 8'b00100000;
		color_arr[7837] = 8'b00100000;
		color_arr[7838] = 8'b00100000;
		color_arr[7839] = 8'b00100000;
		color_arr[7840] = 8'b00100000;
		color_arr[7841] = 8'b00100000;
		color_arr[7842] = 8'b00100000;
		color_arr[7843] = 8'b00100000;
		color_arr[7844] = 8'b00100000;
		color_arr[7845] = 8'b00100000;
		color_arr[7846] = 8'b00100000;
		color_arr[7847] = 8'b00100000;
		color_arr[7848] = 8'b00100000;
		color_arr[7849] = 8'b00100000;
		color_arr[7850] = 8'b00100000;
		color_arr[7851] = 8'b00100000;
		color_arr[7852] = 8'b00100000;
		color_arr[7853] = 8'b00100000;
		color_arr[7854] = 8'b00100000;
		color_arr[7855] = 8'b00100000;
		color_arr[7856] = 8'b00100000;
		color_arr[7857] = 8'b00100000;
		color_arr[7858] = 8'b00100000;
		color_arr[7859] = 8'b00100000;
		color_arr[7860] = 8'b00100000;
		color_arr[7861] = 8'b00100000;
		color_arr[7862] = 8'b00100000;
		color_arr[7863] = 8'b00100000;
		color_arr[7864] = 8'b00100000;
		color_arr[7865] = 8'b00100000;
		color_arr[7866] = 8'b00100000;
		color_arr[7867] = 8'b00100000;
		color_arr[7868] = 8'b00100000;
		color_arr[7869] = 8'b00100000;
		color_arr[7870] = 8'b00100000;
		color_arr[7871] = 8'b00100000;
		color_arr[7872] = 8'b00100000;
		color_arr[7873] = 8'b00100000;
		color_arr[7874] = 8'b00100000;
		color_arr[7875] = 8'b00100000;
		color_arr[7876] = 8'b00100000;
		color_arr[7877] = 8'b00100000;
		color_arr[7878] = 8'b00100000;
		color_arr[7879] = 8'b00100000;
		color_arr[7880] = 8'b00100000;
		color_arr[7881] = 8'b00100000;
		color_arr[7882] = 8'b00100000;
		color_arr[7883] = 8'b00100000;
		color_arr[7884] = 8'b00100000;
		color_arr[7885] = 8'b00100000;
		color_arr[7886] = 8'b00100000;
		color_arr[7887] = 8'b00100000;
		color_arr[7888] = 8'b00001000;
		color_arr[7889] = 8'b00001000;
		color_arr[7890] = 8'b00001000;
		color_arr[7891] = 8'b00001000;
		color_arr[7892] = 8'b00001000;
		color_arr[7893] = 8'b00001000;
		color_arr[7894] = 8'b00001000;
		color_arr[7895] = 8'b00001000;
		color_arr[7896] = 8'b00001000;
		color_arr[7897] = 8'b00001000;
		color_arr[7898] = 8'b00001000;
		color_arr[7899] = 8'b00001000;
		color_arr[7900] = 8'b00001000;
		color_arr[7901] = 8'b00000000;
		color_arr[7902] = 8'b00000000;
		color_arr[7903] = 8'b00001000;
		color_arr[7904] = 8'b00001000;
		color_arr[7905] = 8'b00001000;
		color_arr[7906] = 8'b00001000;
		color_arr[7907] = 8'b00001000;
		color_arr[7908] = 8'b00001000;
		color_arr[7909] = 8'b00001000;
		color_arr[7910] = 8'b00001000;
		color_arr[7911] = 8'b00001000;
		color_arr[7912] = 8'b00001000;
		color_arr[7913] = 8'b00001000;
		color_arr[7914] = 8'b00001000;
		color_arr[7915] = 8'b00001000;
		color_arr[7916] = 8'b00001000;
		color_arr[7917] = 8'b00001000;
		color_arr[7918] = 8'b00001000;
		color_arr[7919] = 8'b00000000;
		color_arr[7920] = 8'b00000000;
		color_arr[7921] = 8'b00001000;
		color_arr[7922] = 8'b00001000;
		color_arr[7923] = 8'b00001000;
		color_arr[7924] = 8'b00001000;
		color_arr[7925] = 8'b00000000;
		color_arr[7926] = 8'b00000000;
		color_arr[7927] = 8'b00001000;
		color_arr[7928] = 8'b00001000;
		color_arr[7929] = 8'b00001000;
		color_arr[7930] = 8'b00001000;
		color_arr[7931] = 8'b00001000;
		color_arr[7932] = 8'b00001000;
		color_arr[7933] = 8'b00010010;
		color_arr[7934] = 8'b00010010;
		color_arr[7935] = 8'b00010010;
		color_arr[7936] = 8'b00010010;
		color_arr[7937] = 8'b00010010;
		color_arr[7938] = 8'b00000000;
		color_arr[7939] = 8'b00000000;
		color_arr[7940] = 8'b00010010;
		color_arr[7941] = 8'b00010010;
		color_arr[7942] = 8'b00010010;
		color_arr[7943] = 8'b00010010;
		color_arr[7944] = 8'b00010010;
		color_arr[7945] = 8'b00010010;
		color_arr[7946] = 8'b00010010;
		color_arr[7947] = 8'b00010010;
		color_arr[7948] = 8'b00010010;
		color_arr[7949] = 8'b00010010;
		color_arr[7950] = 8'b00010010;
		color_arr[7951] = 8'b00010010;
		color_arr[7952] = 8'b00010010;
		color_arr[7953] = 8'b00010010;
		color_arr[7954] = 8'b00100000;
		color_arr[7955] = 8'b00100000;
		color_arr[7956] = 8'b00100000;
		color_arr[7957] = 8'b00000000;
		color_arr[7958] = 8'b00000000;
		color_arr[7959] = 8'b00100000;
		color_arr[7960] = 8'b00100000;
		color_arr[7961] = 8'b00100000;
		color_arr[7962] = 8'b00100000;
		color_arr[7963] = 8'b00100000;
		color_arr[7964] = 8'b00100000;
		color_arr[7965] = 8'b00100000;
		color_arr[7966] = 8'b00100000;
		color_arr[7967] = 8'b00100000;
		color_arr[7968] = 8'b00100000;
		color_arr[7969] = 8'b00100000;
		color_arr[7970] = 8'b00100000;
		color_arr[7971] = 8'b00100000;
		color_arr[7972] = 8'b00100000;
		color_arr[7973] = 8'b00100000;
		color_arr[7974] = 8'b00100000;
		color_arr[7975] = 8'b00100000;
		color_arr[7976] = 8'b00100000;
		color_arr[7977] = 8'b00100000;
		color_arr[7978] = 8'b00100000;
		color_arr[7979] = 8'b00100000;
		color_arr[7980] = 8'b00100000;
		color_arr[7981] = 8'b00100000;
		color_arr[7982] = 8'b00100000;
		color_arr[7983] = 8'b00100000;
		color_arr[7984] = 8'b00100000;
		color_arr[7985] = 8'b00100000;
		color_arr[7986] = 8'b00100000;
		color_arr[7987] = 8'b00100000;
		color_arr[7988] = 8'b00100000;
		color_arr[7989] = 8'b00100000;
		color_arr[7990] = 8'b00100000;
		color_arr[7991] = 8'b00100000;
		color_arr[7992] = 8'b00100000;
		color_arr[7993] = 8'b00100000;
		color_arr[7994] = 8'b00100000;
		color_arr[7995] = 8'b00100000;
		color_arr[7996] = 8'b00100000;
		color_arr[7997] = 8'b00100000;
		color_arr[7998] = 8'b00100000;
		color_arr[7999] = 8'b00100000;
		color_arr[8000] = 8'b00100000;
		color_arr[8001] = 8'b00100000;
		color_arr[8002] = 8'b00100000;
		color_arr[8003] = 8'b00100000;
		color_arr[8004] = 8'b00100000;
		color_arr[8005] = 8'b00100000;
		color_arr[8006] = 8'b00100000;
		color_arr[8007] = 8'b00100000;
		color_arr[8008] = 8'b00100000;
		color_arr[8009] = 8'b00100000;
		color_arr[8010] = 8'b00100000;
		color_arr[8011] = 8'b00100000;
		color_arr[8012] = 8'b00100000;
		color_arr[8013] = 8'b00100000;
		color_arr[8014] = 8'b00100000;
		color_arr[8015] = 8'b00100000;
		color_arr[8016] = 8'b00001000;
		color_arr[8017] = 8'b00001000;
		color_arr[8018] = 8'b00001000;
		color_arr[8019] = 8'b00001000;
		color_arr[8020] = 8'b00001000;
		color_arr[8021] = 8'b00001000;
		color_arr[8022] = 8'b00001000;
		color_arr[8023] = 8'b00001000;
		color_arr[8024] = 8'b00001000;
		color_arr[8025] = 8'b00001000;
		color_arr[8026] = 8'b00001000;
		color_arr[8027] = 8'b00001000;
		color_arr[8028] = 8'b00000000;
		color_arr[8029] = 8'b00000000;
		color_arr[8030] = 8'b00000000;
		color_arr[8031] = 8'b00001000;
		color_arr[8032] = 8'b00001000;
		color_arr[8033] = 8'b00001000;
		color_arr[8034] = 8'b00001000;
		color_arr[8035] = 8'b00001000;
		color_arr[8036] = 8'b00001000;
		color_arr[8037] = 8'b00001000;
		color_arr[8038] = 8'b00001000;
		color_arr[8039] = 8'b00001000;
		color_arr[8040] = 8'b00001000;
		color_arr[8041] = 8'b00001000;
		color_arr[8042] = 8'b00001000;
		color_arr[8043] = 8'b00001000;
		color_arr[8044] = 8'b00001000;
		color_arr[8045] = 8'b00001000;
		color_arr[8046] = 8'b00001000;
		color_arr[8047] = 8'b00000000;
		color_arr[8048] = 8'b00000000;
		color_arr[8049] = 8'b00000000;
		color_arr[8050] = 8'b00001000;
		color_arr[8051] = 8'b00001000;
		color_arr[8052] = 8'b00001000;
		color_arr[8053] = 8'b00000000;
		color_arr[8054] = 8'b00000000;
		color_arr[8055] = 8'b00001000;
		color_arr[8056] = 8'b00001000;
		color_arr[8057] = 8'b00001000;
		color_arr[8058] = 8'b00001000;
		color_arr[8059] = 8'b00001000;
		color_arr[8060] = 8'b00001000;
		color_arr[8061] = 8'b00010010;
		color_arr[8062] = 8'b00010010;
		color_arr[8063] = 8'b00010010;
		color_arr[8064] = 8'b00010010;
		color_arr[8065] = 8'b00010010;
		color_arr[8066] = 8'b00000000;
		color_arr[8067] = 8'b00000000;
		color_arr[8068] = 8'b00010010;
		color_arr[8069] = 8'b00010010;
		color_arr[8070] = 8'b00010010;
		color_arr[8071] = 8'b00010010;
		color_arr[8072] = 8'b00010010;
		color_arr[8073] = 8'b00010010;
		color_arr[8074] = 8'b00010010;
		color_arr[8075] = 8'b00010010;
		color_arr[8076] = 8'b00010010;
		color_arr[8077] = 8'b00010010;
		color_arr[8078] = 8'b00010010;
		color_arr[8079] = 8'b00010010;
		color_arr[8080] = 8'b00010010;
		color_arr[8081] = 8'b00010010;
		color_arr[8082] = 8'b00100000;
		color_arr[8083] = 8'b00100000;
		color_arr[8084] = 8'b00100000;
		color_arr[8085] = 8'b00000000;
		color_arr[8086] = 8'b00000000;
		color_arr[8087] = 8'b00100000;
		color_arr[8088] = 8'b00100000;
		color_arr[8089] = 8'b00100000;
		color_arr[8090] = 8'b00100000;
		color_arr[8091] = 8'b00100000;
		color_arr[8092] = 8'b00100000;
		color_arr[8093] = 8'b00100000;
		color_arr[8094] = 8'b00100000;
		color_arr[8095] = 8'b00100000;
		color_arr[8096] = 8'b00100000;
		color_arr[8097] = 8'b00100000;
		color_arr[8098] = 8'b00100000;
		color_arr[8099] = 8'b00100000;
		color_arr[8100] = 8'b00100000;
		color_arr[8101] = 8'b00100000;
		color_arr[8102] = 8'b00100000;
		color_arr[8103] = 8'b00100000;
		color_arr[8104] = 8'b00100000;
		color_arr[8105] = 8'b00100000;
		color_arr[8106] = 8'b00100000;
		color_arr[8107] = 8'b00100000;
		color_arr[8108] = 8'b00100000;
		color_arr[8109] = 8'b00100000;
		color_arr[8110] = 8'b00100000;
		color_arr[8111] = 8'b00100000;
		color_arr[8112] = 8'b00100000;
		color_arr[8113] = 8'b00100000;
		color_arr[8114] = 8'b00100000;
		color_arr[8115] = 8'b00100000;
		color_arr[8116] = 8'b00100000;
		color_arr[8117] = 8'b00100000;
		color_arr[8118] = 8'b00100000;
		color_arr[8119] = 8'b00100000;
		color_arr[8120] = 8'b00100000;
		color_arr[8121] = 8'b00100000;
		color_arr[8122] = 8'b00100000;
		color_arr[8123] = 8'b00100000;
		color_arr[8124] = 8'b00100000;
		color_arr[8125] = 8'b00100000;
		color_arr[8126] = 8'b00100000;
		color_arr[8127] = 8'b00100000;
		color_arr[8128] = 8'b00100000;
		color_arr[8129] = 8'b00100000;
		color_arr[8130] = 8'b00100000;
		color_arr[8131] = 8'b00100000;
		color_arr[8132] = 8'b00100000;
		color_arr[8133] = 8'b00100000;
		color_arr[8134] = 8'b00100000;
		color_arr[8135] = 8'b00100000;
		color_arr[8136] = 8'b00100000;
		color_arr[8137] = 8'b00100000;
		color_arr[8138] = 8'b00100000;
		color_arr[8139] = 8'b00100000;
		color_arr[8140] = 8'b00100000;
		color_arr[8141] = 8'b00100000;
		color_arr[8142] = 8'b00100000;
		color_arr[8143] = 8'b00100000;
		color_arr[8144] = 8'b00001000;
		color_arr[8145] = 8'b00001000;
		color_arr[8146] = 8'b00001000;
		color_arr[8147] = 8'b00001000;
		color_arr[8148] = 8'b00001000;
		color_arr[8149] = 8'b00001000;
		color_arr[8150] = 8'b00001000;
		color_arr[8151] = 8'b00001000;
		color_arr[8152] = 8'b00001000;
		color_arr[8153] = 8'b00001000;
		color_arr[8154] = 8'b00001000;
		color_arr[8155] = 8'b00001000;
		color_arr[8156] = 8'b00000000;
		color_arr[8157] = 8'b00000000;
		color_arr[8158] = 8'b00001000;
		color_arr[8159] = 8'b00001000;
		color_arr[8160] = 8'b00001000;
		color_arr[8161] = 8'b00001000;
		color_arr[8162] = 8'b00001000;
		color_arr[8163] = 8'b00001000;
		color_arr[8164] = 8'b00001000;
		color_arr[8165] = 8'b00001000;
		color_arr[8166] = 8'b00001000;
		color_arr[8167] = 8'b00001000;
		color_arr[8168] = 8'b00001000;
		color_arr[8169] = 8'b00001000;
		color_arr[8170] = 8'b00001000;
		color_arr[8171] = 8'b00001000;
		color_arr[8172] = 8'b00001000;
		color_arr[8173] = 8'b00001000;
		color_arr[8174] = 8'b00001000;
		color_arr[8175] = 8'b00001000;
		color_arr[8176] = 8'b00000000;
		color_arr[8177] = 8'b00000000;
		color_arr[8178] = 8'b00001000;
		color_arr[8179] = 8'b00001000;
		color_arr[8180] = 8'b00001000;
		color_arr[8181] = 8'b00000000;
		color_arr[8182] = 8'b00000000;
		color_arr[8183] = 8'b00001000;
		color_arr[8184] = 8'b00001000;
		color_arr[8185] = 8'b00001000;
		color_arr[8186] = 8'b00001000;
		color_arr[8187] = 8'b00001000;
		color_arr[8188] = 8'b00001000;
		color_arr[8189] = 8'b00010010;
		color_arr[8190] = 8'b00010010;
		color_arr[8191] = 8'b00010010;
		color_arr[8192] = 8'b00010010;
		color_arr[8193] = 8'b00010010;
		color_arr[8194] = 8'b00000000;
		color_arr[8195] = 8'b00000000;
		color_arr[8196] = 8'b00010010;
		color_arr[8197] = 8'b00010010;
		color_arr[8198] = 8'b00010010;
		color_arr[8199] = 8'b00010010;
		color_arr[8200] = 8'b00010010;
		color_arr[8201] = 8'b00010010;
		color_arr[8202] = 8'b00010010;
		color_arr[8203] = 8'b00010010;
		color_arr[8204] = 8'b00010010;
		color_arr[8205] = 8'b00010010;
		color_arr[8206] = 8'b00010010;
		color_arr[8207] = 8'b00010010;
		color_arr[8208] = 8'b00010010;
		color_arr[8209] = 8'b00010010;
		color_arr[8210] = 8'b00100000;
		color_arr[8211] = 8'b00100000;
		color_arr[8212] = 8'b00100000;
		color_arr[8213] = 8'b00000000;
		color_arr[8214] = 8'b00000000;
		color_arr[8215] = 8'b00100000;
		color_arr[8216] = 8'b00100000;
		color_arr[8217] = 8'b00100000;
		color_arr[8218] = 8'b00100000;
		color_arr[8219] = 8'b00100000;
		color_arr[8220] = 8'b00100000;
		color_arr[8221] = 8'b00100000;
		color_arr[8222] = 8'b00100000;
		color_arr[8223] = 8'b00100000;
		color_arr[8224] = 8'b00100000;
		color_arr[8225] = 8'b00100000;
		color_arr[8226] = 8'b00100000;
		color_arr[8227] = 8'b00100000;
		color_arr[8228] = 8'b00100000;
		color_arr[8229] = 8'b00100000;
		color_arr[8230] = 8'b00100000;
		color_arr[8231] = 8'b00100000;
		color_arr[8232] = 8'b00100000;
		color_arr[8233] = 8'b00100000;
		color_arr[8234] = 8'b00100000;
		color_arr[8235] = 8'b00100000;
		color_arr[8236] = 8'b00100000;
		color_arr[8237] = 8'b00100000;
		color_arr[8238] = 8'b00100000;
		color_arr[8239] = 8'b00100000;
		color_arr[8240] = 8'b00100000;
		color_arr[8241] = 8'b00100000;
		color_arr[8242] = 8'b00100000;
		color_arr[8243] = 8'b00100000;
		color_arr[8244] = 8'b00100000;
		color_arr[8245] = 8'b00100000;
		color_arr[8246] = 8'b00100000;
		color_arr[8247] = 8'b00100000;
		color_arr[8248] = 8'b00100000;
		color_arr[8249] = 8'b00100000;
		color_arr[8250] = 8'b00100000;
		color_arr[8251] = 8'b00100000;
		color_arr[8252] = 8'b00100000;
		color_arr[8253] = 8'b00100000;
		color_arr[8254] = 8'b00100000;
		color_arr[8255] = 8'b00100000;
		color_arr[8256] = 8'b00100000;
		color_arr[8257] = 8'b00100000;
		color_arr[8258] = 8'b00100000;
		color_arr[8259] = 8'b00100000;
		color_arr[8260] = 8'b00100000;
		color_arr[8261] = 8'b00100000;
		color_arr[8262] = 8'b00100000;
		color_arr[8263] = 8'b00100000;
		color_arr[8264] = 8'b00100000;
		color_arr[8265] = 8'b00100000;
		color_arr[8266] = 8'b00100000;
		color_arr[8267] = 8'b00100000;
		color_arr[8268] = 8'b00100000;
		color_arr[8269] = 8'b00100000;
		color_arr[8270] = 8'b00100000;
		color_arr[8271] = 8'b00100000;
		color_arr[8272] = 8'b00001000;
		color_arr[8273] = 8'b00001000;
		color_arr[8274] = 8'b00001000;
		color_arr[8275] = 8'b00001000;
		color_arr[8276] = 8'b00001000;
		color_arr[8277] = 8'b00001000;
		color_arr[8278] = 8'b00001000;
		color_arr[8279] = 8'b00001000;
		color_arr[8280] = 8'b00001000;
		color_arr[8281] = 8'b00001000;
		color_arr[8282] = 8'b00001000;
		color_arr[8283] = 8'b00000000;
		color_arr[8284] = 8'b00000000;
		color_arr[8285] = 8'b00000000;
		color_arr[8286] = 8'b00001000;
		color_arr[8287] = 8'b00001000;
		color_arr[8288] = 8'b00001000;
		color_arr[8289] = 8'b00001000;
		color_arr[8290] = 8'b00001000;
		color_arr[8291] = 8'b00001000;
		color_arr[8292] = 8'b00001000;
		color_arr[8293] = 8'b00001000;
		color_arr[8294] = 8'b00001000;
		color_arr[8295] = 8'b00001000;
		color_arr[8296] = 8'b00001000;
		color_arr[8297] = 8'b00001000;
		color_arr[8298] = 8'b00001000;
		color_arr[8299] = 8'b00001000;
		color_arr[8300] = 8'b00001000;
		color_arr[8301] = 8'b00001000;
		color_arr[8302] = 8'b00001000;
		color_arr[8303] = 8'b00001000;
		color_arr[8304] = 8'b00000000;
		color_arr[8305] = 8'b00000000;
		color_arr[8306] = 8'b00000000;
		color_arr[8307] = 8'b00001000;
		color_arr[8308] = 8'b00001000;
		color_arr[8309] = 8'b00000000;
		color_arr[8310] = 8'b00000000;
		color_arr[8311] = 8'b00001000;
		color_arr[8312] = 8'b00001000;
		color_arr[8313] = 8'b00001000;
		color_arr[8314] = 8'b00001000;
		color_arr[8315] = 8'b00001000;
		color_arr[8316] = 8'b00001000;
		color_arr[8317] = 8'b00010010;
		color_arr[8318] = 8'b00010010;
		color_arr[8319] = 8'b00010010;
		color_arr[8320] = 8'b00010010;
		color_arr[8321] = 8'b00010010;
		color_arr[8322] = 8'b00000000;
		color_arr[8323] = 8'b00000000;
		color_arr[8324] = 8'b00010010;
		color_arr[8325] = 8'b00010010;
		color_arr[8326] = 8'b00010010;
		color_arr[8327] = 8'b00010010;
		color_arr[8328] = 8'b00010010;
		color_arr[8329] = 8'b00010010;
		color_arr[8330] = 8'b00010010;
		color_arr[8331] = 8'b00010010;
		color_arr[8332] = 8'b00010010;
		color_arr[8333] = 8'b00010010;
		color_arr[8334] = 8'b00010010;
		color_arr[8335] = 8'b00010010;
		color_arr[8336] = 8'b00010010;
		color_arr[8337] = 8'b00010010;
		color_arr[8338] = 8'b00100000;
		color_arr[8339] = 8'b00100000;
		color_arr[8340] = 8'b00100000;
		color_arr[8341] = 8'b00000000;
		color_arr[8342] = 8'b00000000;
		color_arr[8343] = 8'b00100000;
		color_arr[8344] = 8'b00100000;
		color_arr[8345] = 8'b00100000;
		color_arr[8346] = 8'b00100000;
		color_arr[8347] = 8'b00100000;
		color_arr[8348] = 8'b00100000;
		color_arr[8349] = 8'b00100000;
		color_arr[8350] = 8'b00100000;
		color_arr[8351] = 8'b00100000;
		color_arr[8352] = 8'b00100000;
		color_arr[8353] = 8'b00100000;
		color_arr[8354] = 8'b00100000;
		color_arr[8355] = 8'b00100000;
		color_arr[8356] = 8'b00100000;
		color_arr[8357] = 8'b00100000;
		color_arr[8358] = 8'b00100000;
		color_arr[8359] = 8'b00100000;
		color_arr[8360] = 8'b00100000;
		color_arr[8361] = 8'b00100000;
		color_arr[8362] = 8'b00100000;
		color_arr[8363] = 8'b00100000;
		color_arr[8364] = 8'b00100000;
		color_arr[8365] = 8'b00100000;
		color_arr[8366] = 8'b00100000;
		color_arr[8367] = 8'b00100000;
		color_arr[8368] = 8'b00100000;
		color_arr[8369] = 8'b00100000;
		color_arr[8370] = 8'b00100000;
		color_arr[8371] = 8'b00100000;
		color_arr[8372] = 8'b00100000;
		color_arr[8373] = 8'b00100000;
		color_arr[8374] = 8'b00100000;
		color_arr[8375] = 8'b00100000;
		color_arr[8376] = 8'b00100000;
		color_arr[8377] = 8'b00100000;
		color_arr[8378] = 8'b00100000;
		color_arr[8379] = 8'b00100000;
		color_arr[8380] = 8'b00100000;
		color_arr[8381] = 8'b00100000;
		color_arr[8382] = 8'b00100000;
		color_arr[8383] = 8'b00100000;
		color_arr[8384] = 8'b00100000;
		color_arr[8385] = 8'b00100000;
		color_arr[8386] = 8'b00100000;
		color_arr[8387] = 8'b00100000;
		color_arr[8388] = 8'b00100000;
		color_arr[8389] = 8'b00100000;
		color_arr[8390] = 8'b00100000;
		color_arr[8391] = 8'b00100000;
		color_arr[8392] = 8'b00100000;
		color_arr[8393] = 8'b00100000;
		color_arr[8394] = 8'b00100000;
		color_arr[8395] = 8'b00100000;
		color_arr[8396] = 8'b00100000;
		color_arr[8397] = 8'b00100000;
		color_arr[8398] = 8'b00100000;
		color_arr[8399] = 8'b00100000;
		color_arr[8400] = 8'b00001000;
		color_arr[8401] = 8'b00001000;
		color_arr[8402] = 8'b00001000;
		color_arr[8403] = 8'b00001000;
		color_arr[8404] = 8'b00001000;
		color_arr[8405] = 8'b00001000;
		color_arr[8406] = 8'b00001000;
		color_arr[8407] = 8'b00001000;
		color_arr[8408] = 8'b00001000;
		color_arr[8409] = 8'b00001000;
		color_arr[8410] = 8'b00000000;
		color_arr[8411] = 8'b00000000;
		color_arr[8412] = 8'b00000000;
		color_arr[8413] = 8'b00001000;
		color_arr[8414] = 8'b00001000;
		color_arr[8415] = 8'b00001000;
		color_arr[8416] = 8'b00001000;
		color_arr[8417] = 8'b00001000;
		color_arr[8418] = 8'b00001000;
		color_arr[8419] = 8'b00001000;
		color_arr[8420] = 8'b00001000;
		color_arr[8421] = 8'b00001000;
		color_arr[8422] = 8'b00001000;
		color_arr[8423] = 8'b00001000;
		color_arr[8424] = 8'b00001000;
		color_arr[8425] = 8'b00001000;
		color_arr[8426] = 8'b00001000;
		color_arr[8427] = 8'b00001000;
		color_arr[8428] = 8'b00001000;
		color_arr[8429] = 8'b00001000;
		color_arr[8430] = 8'b00001000;
		color_arr[8431] = 8'b00001000;
		color_arr[8432] = 8'b00001000;
		color_arr[8433] = 8'b00000000;
		color_arr[8434] = 8'b00000000;
		color_arr[8435] = 8'b00001000;
		color_arr[8436] = 8'b00001000;
		color_arr[8437] = 8'b00000000;
		color_arr[8438] = 8'b00000000;
		color_arr[8439] = 8'b00001000;
		color_arr[8440] = 8'b00001000;
		color_arr[8441] = 8'b00001000;
		color_arr[8442] = 8'b00001000;
		color_arr[8443] = 8'b00001000;
		color_arr[8444] = 8'b00001000;
		color_arr[8445] = 8'b00010010;
		color_arr[8446] = 8'b00010010;
		color_arr[8447] = 8'b00010010;
		color_arr[8448] = 8'b00010010;
		color_arr[8449] = 8'b00010010;
		color_arr[8450] = 8'b00000000;
		color_arr[8451] = 8'b00000000;
		color_arr[8452] = 8'b00010010;
		color_arr[8453] = 8'b00010010;
		color_arr[8454] = 8'b00010010;
		color_arr[8455] = 8'b00010010;
		color_arr[8456] = 8'b00010010;
		color_arr[8457] = 8'b00010010;
		color_arr[8458] = 8'b00010010;
		color_arr[8459] = 8'b00010010;
		color_arr[8460] = 8'b00010010;
		color_arr[8461] = 8'b00010010;
		color_arr[8462] = 8'b00010010;
		color_arr[8463] = 8'b00010010;
		color_arr[8464] = 8'b00010010;
		color_arr[8465] = 8'b00010010;
		color_arr[8466] = 8'b00100000;
		color_arr[8467] = 8'b00100000;
		color_arr[8468] = 8'b00100000;
		color_arr[8469] = 8'b00000000;
		color_arr[8470] = 8'b00000000;
		color_arr[8471] = 8'b00100000;
		color_arr[8472] = 8'b00100000;
		color_arr[8473] = 8'b00100000;
		color_arr[8474] = 8'b00100000;
		color_arr[8475] = 8'b00100000;
		color_arr[8476] = 8'b00100000;
		color_arr[8477] = 8'b00100000;
		color_arr[8478] = 8'b00100000;
		color_arr[8479] = 8'b00100000;
		color_arr[8480] = 8'b00100000;
		color_arr[8481] = 8'b00100000;
		color_arr[8482] = 8'b00100000;
		color_arr[8483] = 8'b00100000;
		color_arr[8484] = 8'b00100000;
		color_arr[8485] = 8'b00100000;
		color_arr[8486] = 8'b00100000;
		color_arr[8487] = 8'b00100000;
		color_arr[8488] = 8'b00100000;
		color_arr[8489] = 8'b00100000;
		color_arr[8490] = 8'b00100000;
		color_arr[8491] = 8'b00100000;
		color_arr[8492] = 8'b00100000;
		color_arr[8493] = 8'b00100000;
		color_arr[8494] = 8'b00100000;
		color_arr[8495] = 8'b00100000;
		color_arr[8496] = 8'b00100000;
		color_arr[8497] = 8'b00100000;
		color_arr[8498] = 8'b00100000;
		color_arr[8499] = 8'b00100000;
		color_arr[8500] = 8'b00100000;
		color_arr[8501] = 8'b00100000;
		color_arr[8502] = 8'b00100000;
		color_arr[8503] = 8'b00100000;
		color_arr[8504] = 8'b00100000;
		color_arr[8505] = 8'b00100000;
		color_arr[8506] = 8'b00100000;
		color_arr[8507] = 8'b00100000;
		color_arr[8508] = 8'b00100000;
		color_arr[8509] = 8'b00100000;
		color_arr[8510] = 8'b00100000;
		color_arr[8511] = 8'b00100000;
		color_arr[8512] = 8'b00100000;
		color_arr[8513] = 8'b00100000;
		color_arr[8514] = 8'b00100000;
		color_arr[8515] = 8'b00100000;
		color_arr[8516] = 8'b00100000;
		color_arr[8517] = 8'b00100000;
		color_arr[8518] = 8'b00100000;
		color_arr[8519] = 8'b00100000;
		color_arr[8520] = 8'b00100000;
		color_arr[8521] = 8'b00100000;
		color_arr[8522] = 8'b00100000;
		color_arr[8523] = 8'b00100000;
		color_arr[8524] = 8'b00100000;
		color_arr[8525] = 8'b00100000;
		color_arr[8526] = 8'b00100000;
		color_arr[8527] = 8'b00100000;
		color_arr[8528] = 8'b00001000;
		color_arr[8529] = 8'b00001000;
		color_arr[8530] = 8'b00001000;
		color_arr[8531] = 8'b00001000;
		color_arr[8532] = 8'b00001000;
		color_arr[8533] = 8'b00001000;
		color_arr[8534] = 8'b00001000;
		color_arr[8535] = 8'b00001000;
		color_arr[8536] = 8'b00001000;
		color_arr[8537] = 8'b00001000;
		color_arr[8538] = 8'b00000000;
		color_arr[8539] = 8'b00000000;
		color_arr[8540] = 8'b00001000;
		color_arr[8541] = 8'b00001000;
		color_arr[8542] = 8'b00001000;
		color_arr[8543] = 8'b00001000;
		color_arr[8544] = 8'b00001000;
		color_arr[8545] = 8'b00001000;
		color_arr[8546] = 8'b00001000;
		color_arr[8547] = 8'b00001000;
		color_arr[8548] = 8'b00001000;
		color_arr[8549] = 8'b00001000;
		color_arr[8550] = 8'b00001000;
		color_arr[8551] = 8'b00001000;
		color_arr[8552] = 8'b00001000;
		color_arr[8553] = 8'b00001000;
		color_arr[8554] = 8'b00001000;
		color_arr[8555] = 8'b00001000;
		color_arr[8556] = 8'b00001000;
		color_arr[8557] = 8'b00001000;
		color_arr[8558] = 8'b00001000;
		color_arr[8559] = 8'b00001000;
		color_arr[8560] = 8'b00001000;
		color_arr[8561] = 8'b00000000;
		color_arr[8562] = 8'b00000000;
		color_arr[8563] = 8'b00001000;
		color_arr[8564] = 8'b00001000;
		color_arr[8565] = 8'b00000000;
		color_arr[8566] = 8'b00000000;
		color_arr[8567] = 8'b00000000;
		color_arr[8568] = 8'b00001000;
		color_arr[8569] = 8'b00001000;
		color_arr[8570] = 8'b00001000;
		color_arr[8571] = 8'b00001000;
		color_arr[8572] = 8'b00001000;
		color_arr[8573] = 8'b00010010;
		color_arr[8574] = 8'b00010010;
		color_arr[8575] = 8'b00010010;
		color_arr[8576] = 8'b00010010;
		color_arr[8577] = 8'b00010010;
		color_arr[8578] = 8'b00000000;
		color_arr[8579] = 8'b00000000;
		color_arr[8580] = 8'b00010010;
		color_arr[8581] = 8'b00010010;
		color_arr[8582] = 8'b00010010;
		color_arr[8583] = 8'b00010010;
		color_arr[8584] = 8'b00010010;
		color_arr[8585] = 8'b00010010;
		color_arr[8586] = 8'b00010010;
		color_arr[8587] = 8'b00010010;
		color_arr[8588] = 8'b00010010;
		color_arr[8589] = 8'b00010010;
		color_arr[8590] = 8'b00010010;
		color_arr[8591] = 8'b00010010;
		color_arr[8592] = 8'b00010010;
		color_arr[8593] = 8'b00010010;
		color_arr[8594] = 8'b00100000;
		color_arr[8595] = 8'b00100000;
		color_arr[8596] = 8'b00100000;
		color_arr[8597] = 8'b00000000;
		color_arr[8598] = 8'b00000000;
		color_arr[8599] = 8'b00100000;
		color_arr[8600] = 8'b00100000;
		color_arr[8601] = 8'b00100000;
		color_arr[8602] = 8'b00100000;
		color_arr[8603] = 8'b00100000;
		color_arr[8604] = 8'b00100000;
		color_arr[8605] = 8'b00100000;
		color_arr[8606] = 8'b00100000;
		color_arr[8607] = 8'b00100000;
		color_arr[8608] = 8'b00100000;
		color_arr[8609] = 8'b00100000;
		color_arr[8610] = 8'b00100000;
		color_arr[8611] = 8'b00100000;
		color_arr[8612] = 8'b00100000;
		color_arr[8613] = 8'b00100000;
		color_arr[8614] = 8'b00100000;
		color_arr[8615] = 8'b00100000;
		color_arr[8616] = 8'b00100000;
		color_arr[8617] = 8'b00100000;
		color_arr[8618] = 8'b00100000;
		color_arr[8619] = 8'b00100000;
		color_arr[8620] = 8'b00100000;
		color_arr[8621] = 8'b00100000;
		color_arr[8622] = 8'b00100000;
		color_arr[8623] = 8'b00100000;
		color_arr[8624] = 8'b00100000;
		color_arr[8625] = 8'b00100000;
		color_arr[8626] = 8'b00100000;
		color_arr[8627] = 8'b00100000;
		color_arr[8628] = 8'b00100000;
		color_arr[8629] = 8'b00100000;
		color_arr[8630] = 8'b00100000;
		color_arr[8631] = 8'b00100000;
		color_arr[8632] = 8'b00100000;
		color_arr[8633] = 8'b00100000;
		color_arr[8634] = 8'b00100000;
		color_arr[8635] = 8'b00100000;
		color_arr[8636] = 8'b00100000;
		color_arr[8637] = 8'b00100000;
		color_arr[8638] = 8'b00100000;
		color_arr[8639] = 8'b00100000;
		color_arr[8640] = 8'b00100000;
		color_arr[8641] = 8'b00100000;
		color_arr[8642] = 8'b00100000;
		color_arr[8643] = 8'b00100000;
		color_arr[8644] = 8'b00100000;
		color_arr[8645] = 8'b00100000;
		color_arr[8646] = 8'b00100000;
		color_arr[8647] = 8'b00100000;
		color_arr[8648] = 8'b00100000;
		color_arr[8649] = 8'b00100000;
		color_arr[8650] = 8'b00100000;
		color_arr[8651] = 8'b00100000;
		color_arr[8652] = 8'b00100000;
		color_arr[8653] = 8'b00100000;
		color_arr[8654] = 8'b00100000;
		color_arr[8655] = 8'b00100000;
		color_arr[8656] = 8'b00001000;
		color_arr[8657] = 8'b00001000;
		color_arr[8658] = 8'b00001000;
		color_arr[8659] = 8'b00001000;
		color_arr[8660] = 8'b00001000;
		color_arr[8661] = 8'b00001000;
		color_arr[8662] = 8'b00001000;
		color_arr[8663] = 8'b00001000;
		color_arr[8664] = 8'b00001000;
		color_arr[8665] = 8'b00000000;
		color_arr[8666] = 8'b00000000;
		color_arr[8667] = 8'b00000000;
		color_arr[8668] = 8'b00001000;
		color_arr[8669] = 8'b00001000;
		color_arr[8670] = 8'b00001000;
		color_arr[8671] = 8'b00001000;
		color_arr[8672] = 8'b00001000;
		color_arr[8673] = 8'b00001000;
		color_arr[8674] = 8'b00001000;
		color_arr[8675] = 8'b00001000;
		color_arr[8676] = 8'b00001000;
		color_arr[8677] = 8'b00001000;
		color_arr[8678] = 8'b00001000;
		color_arr[8679] = 8'b00001000;
		color_arr[8680] = 8'b00001000;
		color_arr[8681] = 8'b00001000;
		color_arr[8682] = 8'b00001000;
		color_arr[8683] = 8'b00001000;
		color_arr[8684] = 8'b00001000;
		color_arr[8685] = 8'b00001000;
		color_arr[8686] = 8'b00001000;
		color_arr[8687] = 8'b00001000;
		color_arr[8688] = 8'b00001000;
		color_arr[8689] = 8'b00000000;
		color_arr[8690] = 8'b00000000;
		color_arr[8691] = 8'b00000000;
		color_arr[8692] = 8'b00001000;
		color_arr[8693] = 8'b00001000;
		color_arr[8694] = 8'b00000000;
		color_arr[8695] = 8'b00000000;
		color_arr[8696] = 8'b00001000;
		color_arr[8697] = 8'b00001000;
		color_arr[8698] = 8'b00001000;
		color_arr[8699] = 8'b00001000;
		color_arr[8700] = 8'b00001000;
		color_arr[8701] = 8'b00010010;
		color_arr[8702] = 8'b00010010;
		color_arr[8703] = 8'b00010010;
		color_arr[8704] = 8'b00010010;
		color_arr[8705] = 8'b00010010;
		color_arr[8706] = 8'b00000000;
		color_arr[8707] = 8'b00000000;
		color_arr[8708] = 8'b00010010;
		color_arr[8709] = 8'b00010010;
		color_arr[8710] = 8'b00010010;
		color_arr[8711] = 8'b00010010;
		color_arr[8712] = 8'b00010010;
		color_arr[8713] = 8'b00010010;
		color_arr[8714] = 8'b00010010;
		color_arr[8715] = 8'b00010010;
		color_arr[8716] = 8'b00010010;
		color_arr[8717] = 8'b00010010;
		color_arr[8718] = 8'b00010010;
		color_arr[8719] = 8'b00010010;
		color_arr[8720] = 8'b00010010;
		color_arr[8721] = 8'b00010010;
		color_arr[8722] = 8'b00100000;
		color_arr[8723] = 8'b00100000;
		color_arr[8724] = 8'b00100000;
		color_arr[8725] = 8'b00000000;
		color_arr[8726] = 8'b00000000;
		color_arr[8727] = 8'b00100000;
		color_arr[8728] = 8'b00100000;
		color_arr[8729] = 8'b00100000;
		color_arr[8730] = 8'b00100000;
		color_arr[8731] = 8'b00100000;
		color_arr[8732] = 8'b00100000;
		color_arr[8733] = 8'b00100000;
		color_arr[8734] = 8'b00100000;
		color_arr[8735] = 8'b00100000;
		color_arr[8736] = 8'b00100000;
		color_arr[8737] = 8'b00100000;
		color_arr[8738] = 8'b00100000;
		color_arr[8739] = 8'b00100000;
		color_arr[8740] = 8'b00100000;
		color_arr[8741] = 8'b00100000;
		color_arr[8742] = 8'b00100000;
		color_arr[8743] = 8'b00100000;
		color_arr[8744] = 8'b00100000;
		color_arr[8745] = 8'b00100000;
		color_arr[8746] = 8'b00100000;
		color_arr[8747] = 8'b00100000;
		color_arr[8748] = 8'b00100000;
		color_arr[8749] = 8'b00100000;
		color_arr[8750] = 8'b00100000;
		color_arr[8751] = 8'b00100000;
		color_arr[8752] = 8'b00100000;
		color_arr[8753] = 8'b00100000;
		color_arr[8754] = 8'b00100000;
		color_arr[8755] = 8'b00100000;
		color_arr[8756] = 8'b00100000;
		color_arr[8757] = 8'b00100000;
		color_arr[8758] = 8'b00100000;
		color_arr[8759] = 8'b00100000;
		color_arr[8760] = 8'b00100000;
		color_arr[8761] = 8'b00100000;
		color_arr[8762] = 8'b00100000;
		color_arr[8763] = 8'b00100000;
		color_arr[8764] = 8'b00100000;
		color_arr[8765] = 8'b00100000;
		color_arr[8766] = 8'b00100000;
		color_arr[8767] = 8'b00100000;
		color_arr[8768] = 8'b00100000;
		color_arr[8769] = 8'b00100000;
		color_arr[8770] = 8'b00100000;
		color_arr[8771] = 8'b00100000;
		color_arr[8772] = 8'b00100000;
		color_arr[8773] = 8'b00100000;
		color_arr[8774] = 8'b00100000;
		color_arr[8775] = 8'b00100000;
		color_arr[8776] = 8'b00100000;
		color_arr[8777] = 8'b00100000;
		color_arr[8778] = 8'b00100000;
		color_arr[8779] = 8'b00100000;
		color_arr[8780] = 8'b00100000;
		color_arr[8781] = 8'b00100000;
		color_arr[8782] = 8'b00100000;
		color_arr[8783] = 8'b00100000;
		color_arr[8784] = 8'b00001000;
		color_arr[8785] = 8'b00001000;
		color_arr[8786] = 8'b00001000;
		color_arr[8787] = 8'b00001000;
		color_arr[8788] = 8'b00001000;
		color_arr[8789] = 8'b00001000;
		color_arr[8790] = 8'b00001000;
		color_arr[8791] = 8'b00001000;
		color_arr[8792] = 8'b00001000;
		color_arr[8793] = 8'b00000000;
		color_arr[8794] = 8'b00000000;
		color_arr[8795] = 8'b00001000;
		color_arr[8796] = 8'b00001000;
		color_arr[8797] = 8'b00001000;
		color_arr[8798] = 8'b00001000;
		color_arr[8799] = 8'b00001000;
		color_arr[8800] = 8'b00001000;
		color_arr[8801] = 8'b00001000;
		color_arr[8802] = 8'b00001000;
		color_arr[8803] = 8'b00001000;
		color_arr[8804] = 8'b00001000;
		color_arr[8805] = 8'b00001000;
		color_arr[8806] = 8'b00001000;
		color_arr[8807] = 8'b00001000;
		color_arr[8808] = 8'b00001000;
		color_arr[8809] = 8'b00001000;
		color_arr[8810] = 8'b00001000;
		color_arr[8811] = 8'b00001000;
		color_arr[8812] = 8'b00001000;
		color_arr[8813] = 8'b00001000;
		color_arr[8814] = 8'b00001000;
		color_arr[8815] = 8'b00001000;
		color_arr[8816] = 8'b00001000;
		color_arr[8817] = 8'b00001000;
		color_arr[8818] = 8'b00000000;
		color_arr[8819] = 8'b00000000;
		color_arr[8820] = 8'b00001000;
		color_arr[8821] = 8'b00001000;
		color_arr[8822] = 8'b00000000;
		color_arr[8823] = 8'b00000000;
		color_arr[8824] = 8'b00001000;
		color_arr[8825] = 8'b00001000;
		color_arr[8826] = 8'b00001000;
		color_arr[8827] = 8'b00001000;
		color_arr[8828] = 8'b00001000;
		color_arr[8829] = 8'b00010010;
		color_arr[8830] = 8'b00010010;
		color_arr[8831] = 8'b00010010;
		color_arr[8832] = 8'b00010010;
		color_arr[8833] = 8'b00010010;
		color_arr[8834] = 8'b00000000;
		color_arr[8835] = 8'b00000000;
		color_arr[8836] = 8'b00010010;
		color_arr[8837] = 8'b00010010;
		color_arr[8838] = 8'b00010010;
		color_arr[8839] = 8'b00010010;
		color_arr[8840] = 8'b00010010;
		color_arr[8841] = 8'b00010010;
		color_arr[8842] = 8'b00010010;
		color_arr[8843] = 8'b00010010;
		color_arr[8844] = 8'b00010010;
		color_arr[8845] = 8'b00010010;
		color_arr[8846] = 8'b00010010;
		color_arr[8847] = 8'b00010010;
		color_arr[8848] = 8'b00010010;
		color_arr[8849] = 8'b00010010;
		color_arr[8850] = 8'b00100000;
		color_arr[8851] = 8'b00100000;
		color_arr[8852] = 8'b00100000;
		color_arr[8853] = 8'b00000000;
		color_arr[8854] = 8'b00000000;
		color_arr[8855] = 8'b00100000;
		color_arr[8856] = 8'b00100000;
		color_arr[8857] = 8'b00100000;
		color_arr[8858] = 8'b00100000;
		color_arr[8859] = 8'b00100000;
		color_arr[8860] = 8'b00100000;
		color_arr[8861] = 8'b00100000;
		color_arr[8862] = 8'b00100000;
		color_arr[8863] = 8'b00100000;
		color_arr[8864] = 8'b00100000;
		color_arr[8865] = 8'b00100000;
		color_arr[8866] = 8'b00100000;
		color_arr[8867] = 8'b00100000;
		color_arr[8868] = 8'b00100000;
		color_arr[8869] = 8'b00100000;
		color_arr[8870] = 8'b00100000;
		color_arr[8871] = 8'b00100000;
		color_arr[8872] = 8'b00100000;
		color_arr[8873] = 8'b00100000;
		color_arr[8874] = 8'b00100000;
		color_arr[8875] = 8'b00100000;
		color_arr[8876] = 8'b00100000;
		color_arr[8877] = 8'b00100000;
		color_arr[8878] = 8'b00100000;
		color_arr[8879] = 8'b00100000;
		color_arr[8880] = 8'b00100000;
		color_arr[8881] = 8'b00100000;
		color_arr[8882] = 8'b00100000;
		color_arr[8883] = 8'b00100000;
		color_arr[8884] = 8'b00100000;
		color_arr[8885] = 8'b00100000;
		color_arr[8886] = 8'b00100000;
		color_arr[8887] = 8'b00100000;
		color_arr[8888] = 8'b00100000;
		color_arr[8889] = 8'b00100000;
		color_arr[8890] = 8'b00100000;
		color_arr[8891] = 8'b00100000;
		color_arr[8892] = 8'b00100000;
		color_arr[8893] = 8'b00100000;
		color_arr[8894] = 8'b00100000;
		color_arr[8895] = 8'b00100000;
		color_arr[8896] = 8'b00100000;
		color_arr[8897] = 8'b00100000;
		color_arr[8898] = 8'b00100000;
		color_arr[8899] = 8'b00100000;
		color_arr[8900] = 8'b00100000;
		color_arr[8901] = 8'b00100000;
		color_arr[8902] = 8'b00100000;
		color_arr[8903] = 8'b00100000;
		color_arr[8904] = 8'b00100000;
		color_arr[8905] = 8'b00100000;
		color_arr[8906] = 8'b00100000;
		color_arr[8907] = 8'b00100000;
		color_arr[8908] = 8'b00100000;
		color_arr[8909] = 8'b00100000;
		color_arr[8910] = 8'b00100000;
		color_arr[8911] = 8'b00100000;
		color_arr[8912] = 8'b00001000;
		color_arr[8913] = 8'b00001000;
		color_arr[8914] = 8'b00001000;
		color_arr[8915] = 8'b00001000;
		color_arr[8916] = 8'b00001000;
		color_arr[8917] = 8'b00001000;
		color_arr[8918] = 8'b00001000;
		color_arr[8919] = 8'b00001000;
		color_arr[8920] = 8'b00000000;
		color_arr[8921] = 8'b00000000;
		color_arr[8922] = 8'b00000000;
		color_arr[8923] = 8'b00001000;
		color_arr[8924] = 8'b00001000;
		color_arr[8925] = 8'b00001000;
		color_arr[8926] = 8'b00001000;
		color_arr[8927] = 8'b00001000;
		color_arr[8928] = 8'b00001000;
		color_arr[8929] = 8'b00001000;
		color_arr[8930] = 8'b00001000;
		color_arr[8931] = 8'b00001000;
		color_arr[8932] = 8'b00001000;
		color_arr[8933] = 8'b00001000;
		color_arr[8934] = 8'b00001000;
		color_arr[8935] = 8'b00001000;
		color_arr[8936] = 8'b00001000;
		color_arr[8937] = 8'b00001000;
		color_arr[8938] = 8'b00001000;
		color_arr[8939] = 8'b00001000;
		color_arr[8940] = 8'b00001000;
		color_arr[8941] = 8'b00001000;
		color_arr[8942] = 8'b00001000;
		color_arr[8943] = 8'b00001000;
		color_arr[8944] = 8'b00001000;
		color_arr[8945] = 8'b00001000;
		color_arr[8946] = 8'b00000000;
		color_arr[8947] = 8'b00000000;
		color_arr[8948] = 8'b00000000;
		color_arr[8949] = 8'b00001000;
		color_arr[8950] = 8'b00000000;
		color_arr[8951] = 8'b00000000;
		color_arr[8952] = 8'b00001000;
		color_arr[8953] = 8'b00001000;
		color_arr[8954] = 8'b00001000;
		color_arr[8955] = 8'b00001000;
		color_arr[8956] = 8'b00001000;
		color_arr[8957] = 8'b00010010;
		color_arr[8958] = 8'b00010010;
		color_arr[8959] = 8'b00010010;
		color_arr[8960] = 8'b00010010;
		color_arr[8961] = 8'b00010010;
		color_arr[8962] = 8'b00000000;
		color_arr[8963] = 8'b00000000;
		color_arr[8964] = 8'b00010010;
		color_arr[8965] = 8'b00010010;
		color_arr[8966] = 8'b00010010;
		color_arr[8967] = 8'b00010010;
		color_arr[8968] = 8'b00010010;
		color_arr[8969] = 8'b00010010;
		color_arr[8970] = 8'b00010010;
		color_arr[8971] = 8'b00010010;
		color_arr[8972] = 8'b00010010;
		color_arr[8973] = 8'b00010010;
		color_arr[8974] = 8'b00010010;
		color_arr[8975] = 8'b00010010;
		color_arr[8976] = 8'b00010010;
		color_arr[8977] = 8'b00010010;
		color_arr[8978] = 8'b00100000;
		color_arr[8979] = 8'b00100000;
		color_arr[8980] = 8'b00100000;
		color_arr[8981] = 8'b00000000;
		color_arr[8982] = 8'b00000000;
		color_arr[8983] = 8'b00100000;
		color_arr[8984] = 8'b00100000;
		color_arr[8985] = 8'b00100000;
		color_arr[8986] = 8'b00100000;
		color_arr[8987] = 8'b00100000;
		color_arr[8988] = 8'b00100000;
		color_arr[8989] = 8'b00100000;
		color_arr[8990] = 8'b00100000;
		color_arr[8991] = 8'b00100000;
		color_arr[8992] = 8'b00100000;
		color_arr[8993] = 8'b00100000;
		color_arr[8994] = 8'b00100000;
		color_arr[8995] = 8'b00100000;
		color_arr[8996] = 8'b00100000;
		color_arr[8997] = 8'b00100000;
		color_arr[8998] = 8'b00100000;
		color_arr[8999] = 8'b00100000;
		color_arr[9000] = 8'b00100000;
		color_arr[9001] = 8'b00100000;
		color_arr[9002] = 8'b00100000;
		color_arr[9003] = 8'b00100000;
		color_arr[9004] = 8'b00100000;
		color_arr[9005] = 8'b00100000;
		color_arr[9006] = 8'b00100000;
		color_arr[9007] = 8'b00100000;
		color_arr[9008] = 8'b00100000;
		color_arr[9009] = 8'b00100000;
		color_arr[9010] = 8'b00100000;
		color_arr[9011] = 8'b00100000;
		color_arr[9012] = 8'b00100000;
		color_arr[9013] = 8'b00100000;
		color_arr[9014] = 8'b00100000;
		color_arr[9015] = 8'b00100000;
		color_arr[9016] = 8'b00100000;
		color_arr[9017] = 8'b00100000;
		color_arr[9018] = 8'b00100000;
		color_arr[9019] = 8'b00100000;
		color_arr[9020] = 8'b00100000;
		color_arr[9021] = 8'b00100000;
		color_arr[9022] = 8'b00100000;
		color_arr[9023] = 8'b00100000;
		color_arr[9024] = 8'b00100000;
		color_arr[9025] = 8'b00100000;
		color_arr[9026] = 8'b00100000;
		color_arr[9027] = 8'b00100000;
		color_arr[9028] = 8'b00100000;
		color_arr[9029] = 8'b00100000;
		color_arr[9030] = 8'b00100000;
		color_arr[9031] = 8'b00100000;
		color_arr[9032] = 8'b00100000;
		color_arr[9033] = 8'b00100000;
		color_arr[9034] = 8'b00100000;
		color_arr[9035] = 8'b00100000;
		color_arr[9036] = 8'b00100000;
		color_arr[9037] = 8'b00100000;
		color_arr[9038] = 8'b00100000;
		color_arr[9039] = 8'b00100000;
		color_arr[9040] = 8'b00001000;
		color_arr[9041] = 8'b00001000;
		color_arr[9042] = 8'b00001000;
		color_arr[9043] = 8'b00001000;
		color_arr[9044] = 8'b00001000;
		color_arr[9045] = 8'b00001000;
		color_arr[9046] = 8'b00001000;
		color_arr[9047] = 8'b00001000;
		color_arr[9048] = 8'b00000000;
		color_arr[9049] = 8'b00000000;
		color_arr[9050] = 8'b00001000;
		color_arr[9051] = 8'b00001000;
		color_arr[9052] = 8'b00001000;
		color_arr[9053] = 8'b00001000;
		color_arr[9054] = 8'b00001000;
		color_arr[9055] = 8'b00001000;
		color_arr[9056] = 8'b00001000;
		color_arr[9057] = 8'b00001000;
		color_arr[9058] = 8'b00001000;
		color_arr[9059] = 8'b00001000;
		color_arr[9060] = 8'b00001000;
		color_arr[9061] = 8'b00001000;
		color_arr[9062] = 8'b00001000;
		color_arr[9063] = 8'b00001000;
		color_arr[9064] = 8'b00001000;
		color_arr[9065] = 8'b00001000;
		color_arr[9066] = 8'b00001000;
		color_arr[9067] = 8'b00001000;
		color_arr[9068] = 8'b00001000;
		color_arr[9069] = 8'b00001000;
		color_arr[9070] = 8'b00001000;
		color_arr[9071] = 8'b00001000;
		color_arr[9072] = 8'b00001000;
		color_arr[9073] = 8'b00001000;
		color_arr[9074] = 8'b00001000;
		color_arr[9075] = 8'b00000000;
		color_arr[9076] = 8'b00000000;
		color_arr[9077] = 8'b00001000;
		color_arr[9078] = 8'b00000000;
		color_arr[9079] = 8'b00000000;
		color_arr[9080] = 8'b00001000;
		color_arr[9081] = 8'b00001000;
		color_arr[9082] = 8'b00001000;
		color_arr[9083] = 8'b00001000;
		color_arr[9084] = 8'b00001000;
		color_arr[9085] = 8'b00010010;
		color_arr[9086] = 8'b00010010;
		color_arr[9087] = 8'b00010010;
		color_arr[9088] = 8'b00010010;
		color_arr[9089] = 8'b00010010;
		color_arr[9090] = 8'b00000000;
		color_arr[9091] = 8'b00000000;
		color_arr[9092] = 8'b00010010;
		color_arr[9093] = 8'b00010010;
		color_arr[9094] = 8'b00010010;
		color_arr[9095] = 8'b00010010;
		color_arr[9096] = 8'b00010010;
		color_arr[9097] = 8'b00010010;
		color_arr[9098] = 8'b00010010;
		color_arr[9099] = 8'b00010010;
		color_arr[9100] = 8'b00010010;
		color_arr[9101] = 8'b00010010;
		color_arr[9102] = 8'b00010010;
		color_arr[9103] = 8'b00010010;
		color_arr[9104] = 8'b00010010;
		color_arr[9105] = 8'b00010010;
		color_arr[9106] = 8'b00100000;
		color_arr[9107] = 8'b00100000;
		color_arr[9108] = 8'b00100000;
		color_arr[9109] = 8'b00000000;
		color_arr[9110] = 8'b00000000;
		color_arr[9111] = 8'b00100000;
		color_arr[9112] = 8'b00100000;
		color_arr[9113] = 8'b00100000;
		color_arr[9114] = 8'b00100000;
		color_arr[9115] = 8'b00100000;
		color_arr[9116] = 8'b00100000;
		color_arr[9117] = 8'b00100000;
		color_arr[9118] = 8'b00100000;
		color_arr[9119] = 8'b00100000;
		color_arr[9120] = 8'b00100000;
		color_arr[9121] = 8'b00100000;
		color_arr[9122] = 8'b00100000;
		color_arr[9123] = 8'b00100000;
		color_arr[9124] = 8'b00100000;
		color_arr[9125] = 8'b00100000;
		color_arr[9126] = 8'b00100000;
		color_arr[9127] = 8'b00100000;
		color_arr[9128] = 8'b00100000;
		color_arr[9129] = 8'b00100000;
		color_arr[9130] = 8'b00100000;
		color_arr[9131] = 8'b00100000;
		color_arr[9132] = 8'b00100000;
		color_arr[9133] = 8'b00100000;
		color_arr[9134] = 8'b00100000;
		color_arr[9135] = 8'b00100000;
		color_arr[9136] = 8'b00100000;
		color_arr[9137] = 8'b00100000;
		color_arr[9138] = 8'b00100000;
		color_arr[9139] = 8'b00100000;
		color_arr[9140] = 8'b00100000;
		color_arr[9141] = 8'b00100000;
		color_arr[9142] = 8'b00100000;
		color_arr[9143] = 8'b00100000;
		color_arr[9144] = 8'b00100000;
		color_arr[9145] = 8'b00100000;
		color_arr[9146] = 8'b00100000;
		color_arr[9147] = 8'b00100000;
		color_arr[9148] = 8'b00100000;
		color_arr[9149] = 8'b00100000;
		color_arr[9150] = 8'b00100000;
		color_arr[9151] = 8'b00100000;
		color_arr[9152] = 8'b00100000;
		color_arr[9153] = 8'b00100000;
		color_arr[9154] = 8'b00100000;
		color_arr[9155] = 8'b00100000;
		color_arr[9156] = 8'b00100000;
		color_arr[9157] = 8'b00100000;
		color_arr[9158] = 8'b00100000;
		color_arr[9159] = 8'b00100000;
		color_arr[9160] = 8'b00100000;
		color_arr[9161] = 8'b00100000;
		color_arr[9162] = 8'b00100000;
		color_arr[9163] = 8'b00100000;
		color_arr[9164] = 8'b00100000;
		color_arr[9165] = 8'b00100000;
		color_arr[9166] = 8'b00100000;
		color_arr[9167] = 8'b00100000;
		color_arr[9168] = 8'b00001000;
		color_arr[9169] = 8'b00001000;
		color_arr[9170] = 8'b00001000;
		color_arr[9171] = 8'b00001000;
		color_arr[9172] = 8'b00001000;
		color_arr[9173] = 8'b00001000;
		color_arr[9174] = 8'b00001000;
		color_arr[9175] = 8'b00000000;
		color_arr[9176] = 8'b00000000;
		color_arr[9177] = 8'b00000000;
		color_arr[9178] = 8'b00001000;
		color_arr[9179] = 8'b00001000;
		color_arr[9180] = 8'b00001000;
		color_arr[9181] = 8'b00001000;
		color_arr[9182] = 8'b00001000;
		color_arr[9183] = 8'b00001000;
		color_arr[9184] = 8'b00001000;
		color_arr[9185] = 8'b00001000;
		color_arr[9186] = 8'b00001000;
		color_arr[9187] = 8'b00001000;
		color_arr[9188] = 8'b00001000;
		color_arr[9189] = 8'b00001000;
		color_arr[9190] = 8'b00001000;
		color_arr[9191] = 8'b00001000;
		color_arr[9192] = 8'b00001000;
		color_arr[9193] = 8'b00001000;
		color_arr[9194] = 8'b00001000;
		color_arr[9195] = 8'b00001000;
		color_arr[9196] = 8'b00001000;
		color_arr[9197] = 8'b00001000;
		color_arr[9198] = 8'b00001000;
		color_arr[9199] = 8'b00001000;
		color_arr[9200] = 8'b00001000;
		color_arr[9201] = 8'b00001000;
		color_arr[9202] = 8'b00001000;
		color_arr[9203] = 8'b00000000;
		color_arr[9204] = 8'b00000000;
		color_arr[9205] = 8'b00000000;
		color_arr[9206] = 8'b00000000;
		color_arr[9207] = 8'b00000000;
		color_arr[9208] = 8'b00001000;
		color_arr[9209] = 8'b00001000;
		color_arr[9210] = 8'b00001000;
		color_arr[9211] = 8'b00001000;
		color_arr[9212] = 8'b00001000;
		color_arr[9213] = 8'b00010010;
		color_arr[9214] = 8'b00010010;
		color_arr[9215] = 8'b00010010;
		color_arr[9216] = 8'b00010010;
		color_arr[9217] = 8'b00010010;
		color_arr[9218] = 8'b00000000;
		color_arr[9219] = 8'b00000000;
		color_arr[9220] = 8'b00010010;
		color_arr[9221] = 8'b00010010;
		color_arr[9222] = 8'b00010010;
		color_arr[9223] = 8'b00010010;
		color_arr[9224] = 8'b00010010;
		color_arr[9225] = 8'b00010010;
		color_arr[9226] = 8'b00010010;
		color_arr[9227] = 8'b00010010;
		color_arr[9228] = 8'b00010010;
		color_arr[9229] = 8'b00010010;
		color_arr[9230] = 8'b00010010;
		color_arr[9231] = 8'b00010010;
		color_arr[9232] = 8'b00010010;
		color_arr[9233] = 8'b00010010;
		color_arr[9234] = 8'b00100000;
		color_arr[9235] = 8'b00100000;
		color_arr[9236] = 8'b00100000;
		color_arr[9237] = 8'b00000000;
		color_arr[9238] = 8'b00000000;
		color_arr[9239] = 8'b00100000;
		color_arr[9240] = 8'b00100000;
		color_arr[9241] = 8'b00100000;
		color_arr[9242] = 8'b00100000;
		color_arr[9243] = 8'b00100000;
		color_arr[9244] = 8'b00100000;
		color_arr[9245] = 8'b00100000;
		color_arr[9246] = 8'b00100000;
		color_arr[9247] = 8'b00100000;
		color_arr[9248] = 8'b00100000;
		color_arr[9249] = 8'b00100000;
		color_arr[9250] = 8'b00100000;
		color_arr[9251] = 8'b00100000;
		color_arr[9252] = 8'b00100000;
		color_arr[9253] = 8'b00100000;
		color_arr[9254] = 8'b00100000;
		color_arr[9255] = 8'b00100000;
		color_arr[9256] = 8'b00100000;
		color_arr[9257] = 8'b00100000;
		color_arr[9258] = 8'b00100000;
		color_arr[9259] = 8'b00100000;
		color_arr[9260] = 8'b00100000;
		color_arr[9261] = 8'b00100000;
		color_arr[9262] = 8'b00100000;
		color_arr[9263] = 8'b00100000;
		color_arr[9264] = 8'b00100000;
		color_arr[9265] = 8'b00100000;
		color_arr[9266] = 8'b00100000;
		color_arr[9267] = 8'b00100000;
		color_arr[9268] = 8'b00100000;
		color_arr[9269] = 8'b00100000;
		color_arr[9270] = 8'b00100000;
		color_arr[9271] = 8'b00100000;
		color_arr[9272] = 8'b00100000;
		color_arr[9273] = 8'b00100000;
		color_arr[9274] = 8'b00100000;
		color_arr[9275] = 8'b00100000;
		color_arr[9276] = 8'b00100000;
		color_arr[9277] = 8'b00100000;
		color_arr[9278] = 8'b00100000;
		color_arr[9279] = 8'b00100000;
		color_arr[9280] = 8'b00100000;
		color_arr[9281] = 8'b00100000;
		color_arr[9282] = 8'b00100000;
		color_arr[9283] = 8'b00100000;
		color_arr[9284] = 8'b00100000;
		color_arr[9285] = 8'b00100000;
		color_arr[9286] = 8'b00100000;
		color_arr[9287] = 8'b00100000;
		color_arr[9288] = 8'b00100000;
		color_arr[9289] = 8'b00100000;
		color_arr[9290] = 8'b00100000;
		color_arr[9291] = 8'b00100000;
		color_arr[9292] = 8'b00100000;
		color_arr[9293] = 8'b00100000;
		color_arr[9294] = 8'b00100000;
		color_arr[9295] = 8'b00100000;
		color_arr[9296] = 8'b00001000;
		color_arr[9297] = 8'b00001000;
		color_arr[9298] = 8'b00001000;
		color_arr[9299] = 8'b00001000;
		color_arr[9300] = 8'b00001000;
		color_arr[9301] = 8'b00001000;
		color_arr[9302] = 8'b00000000;
		color_arr[9303] = 8'b00000000;
		color_arr[9304] = 8'b00000000;
		color_arr[9305] = 8'b00001000;
		color_arr[9306] = 8'b00001000;
		color_arr[9307] = 8'b00001000;
		color_arr[9308] = 8'b00001000;
		color_arr[9309] = 8'b00001000;
		color_arr[9310] = 8'b00001000;
		color_arr[9311] = 8'b00001000;
		color_arr[9312] = 8'b00001000;
		color_arr[9313] = 8'b00001000;
		color_arr[9314] = 8'b00001000;
		color_arr[9315] = 8'b00001000;
		color_arr[9316] = 8'b00001000;
		color_arr[9317] = 8'b00001000;
		color_arr[9318] = 8'b00001000;
		color_arr[9319] = 8'b00001000;
		color_arr[9320] = 8'b00001000;
		color_arr[9321] = 8'b00001000;
		color_arr[9322] = 8'b00001000;
		color_arr[9323] = 8'b00001000;
		color_arr[9324] = 8'b00001000;
		color_arr[9325] = 8'b00001000;
		color_arr[9326] = 8'b00001000;
		color_arr[9327] = 8'b00001000;
		color_arr[9328] = 8'b00001000;
		color_arr[9329] = 8'b00001000;
		color_arr[9330] = 8'b00001000;
		color_arr[9331] = 8'b00001000;
		color_arr[9332] = 8'b00000000;
		color_arr[9333] = 8'b00000000;
		color_arr[9334] = 8'b00000000;
		color_arr[9335] = 8'b00000000;
		color_arr[9336] = 8'b00001000;
		color_arr[9337] = 8'b00001000;
		color_arr[9338] = 8'b00001000;
		color_arr[9339] = 8'b00001000;
		color_arr[9340] = 8'b00001000;
		color_arr[9341] = 8'b00010010;
		color_arr[9342] = 8'b00010010;
		color_arr[9343] = 8'b00010010;
		color_arr[9344] = 8'b00010010;
		color_arr[9345] = 8'b00010010;
		color_arr[9346] = 8'b00000000;
		color_arr[9347] = 8'b00000000;
		color_arr[9348] = 8'b00010010;
		color_arr[9349] = 8'b00010010;
		color_arr[9350] = 8'b00010010;
		color_arr[9351] = 8'b00010010;
		color_arr[9352] = 8'b00010010;
		color_arr[9353] = 8'b00010010;
		color_arr[9354] = 8'b00010010;
		color_arr[9355] = 8'b00010010;
		color_arr[9356] = 8'b00010010;
		color_arr[9357] = 8'b00010010;
		color_arr[9358] = 8'b00010010;
		color_arr[9359] = 8'b00010010;
		color_arr[9360] = 8'b00010010;
		color_arr[9361] = 8'b00010010;
		color_arr[9362] = 8'b00100000;
		color_arr[9363] = 8'b00100000;
		color_arr[9364] = 8'b00100000;
		color_arr[9365] = 8'b00000000;
		color_arr[9366] = 8'b00000000;
		color_arr[9367] = 8'b00100000;
		color_arr[9368] = 8'b00100000;
		color_arr[9369] = 8'b00100000;
		color_arr[9370] = 8'b00100000;
		color_arr[9371] = 8'b00100000;
		color_arr[9372] = 8'b00100000;
		color_arr[9373] = 8'b00100000;
		color_arr[9374] = 8'b00100000;
		color_arr[9375] = 8'b00100000;
		color_arr[9376] = 8'b00100000;
		color_arr[9377] = 8'b00100000;
		color_arr[9378] = 8'b00100000;
		color_arr[9379] = 8'b00100000;
		color_arr[9380] = 8'b00100000;
		color_arr[9381] = 8'b00100000;
		color_arr[9382] = 8'b00100000;
		color_arr[9383] = 8'b00100000;
		color_arr[9384] = 8'b00100000;
		color_arr[9385] = 8'b00100000;
		color_arr[9386] = 8'b00100000;
		color_arr[9387] = 8'b00100000;
		color_arr[9388] = 8'b00100000;
		color_arr[9389] = 8'b00100000;
		color_arr[9390] = 8'b00100000;
		color_arr[9391] = 8'b00100000;
		color_arr[9392] = 8'b00100000;
		color_arr[9393] = 8'b00100000;
		color_arr[9394] = 8'b00100000;
		color_arr[9395] = 8'b00100000;
		color_arr[9396] = 8'b00100000;
		color_arr[9397] = 8'b00100000;
		color_arr[9398] = 8'b00100000;
		color_arr[9399] = 8'b00100000;
		color_arr[9400] = 8'b00100000;
		color_arr[9401] = 8'b00100000;
		color_arr[9402] = 8'b00100000;
		color_arr[9403] = 8'b00100000;
		color_arr[9404] = 8'b00100000;
		color_arr[9405] = 8'b00100000;
		color_arr[9406] = 8'b00100000;
		color_arr[9407] = 8'b00100000;
		color_arr[9408] = 8'b00100000;
		color_arr[9409] = 8'b00100000;
		color_arr[9410] = 8'b00100000;
		color_arr[9411] = 8'b00100000;
		color_arr[9412] = 8'b00100000;
		color_arr[9413] = 8'b00100000;
		color_arr[9414] = 8'b00100000;
		color_arr[9415] = 8'b00100000;
		color_arr[9416] = 8'b00100000;
		color_arr[9417] = 8'b00100000;
		color_arr[9418] = 8'b00100000;
		color_arr[9419] = 8'b00100000;
		color_arr[9420] = 8'b00100000;
		color_arr[9421] = 8'b00100000;
		color_arr[9422] = 8'b00100000;
		color_arr[9423] = 8'b00100000;
		color_arr[9424] = 8'b00001000;
		color_arr[9425] = 8'b00001000;
		color_arr[9426] = 8'b00001000;
		color_arr[9427] = 8'b00001000;
		color_arr[9428] = 8'b00001000;
		color_arr[9429] = 8'b00000000;
		color_arr[9430] = 8'b00000000;
		color_arr[9431] = 8'b00000000;
		color_arr[9432] = 8'b00001000;
		color_arr[9433] = 8'b00001000;
		color_arr[9434] = 8'b00001000;
		color_arr[9435] = 8'b00001000;
		color_arr[9436] = 8'b00001000;
		color_arr[9437] = 8'b00001000;
		color_arr[9438] = 8'b00001000;
		color_arr[9439] = 8'b00001000;
		color_arr[9440] = 8'b00001000;
		color_arr[9441] = 8'b00001000;
		color_arr[9442] = 8'b00001000;
		color_arr[9443] = 8'b00001000;
		color_arr[9444] = 8'b00001000;
		color_arr[9445] = 8'b00001000;
		color_arr[9446] = 8'b00001000;
		color_arr[9447] = 8'b00001000;
		color_arr[9448] = 8'b00001000;
		color_arr[9449] = 8'b00001000;
		color_arr[9450] = 8'b00001000;
		color_arr[9451] = 8'b00001000;
		color_arr[9452] = 8'b00001000;
		color_arr[9453] = 8'b00001000;
		color_arr[9454] = 8'b00001000;
		color_arr[9455] = 8'b00001000;
		color_arr[9456] = 8'b00001000;
		color_arr[9457] = 8'b00001000;
		color_arr[9458] = 8'b00001000;
		color_arr[9459] = 8'b00001000;
		color_arr[9460] = 8'b00000000;
		color_arr[9461] = 8'b00000000;
		color_arr[9462] = 8'b00000000;
		color_arr[9463] = 8'b00000000;
		color_arr[9464] = 8'b00000000;
		color_arr[9465] = 8'b00001000;
		color_arr[9466] = 8'b00001000;
		color_arr[9467] = 8'b00001000;
		color_arr[9468] = 8'b00001000;
		color_arr[9469] = 8'b00010010;
		color_arr[9470] = 8'b00010010;
		color_arr[9471] = 8'b00010010;
		color_arr[9472] = 8'b00010010;
		color_arr[9473] = 8'b00010010;
		color_arr[9474] = 8'b00000000;
		color_arr[9475] = 8'b00000000;
		color_arr[9476] = 8'b00010010;
		color_arr[9477] = 8'b00010010;
		color_arr[9478] = 8'b00010010;
		color_arr[9479] = 8'b00010010;
		color_arr[9480] = 8'b00010010;
		color_arr[9481] = 8'b00010010;
		color_arr[9482] = 8'b00010010;
		color_arr[9483] = 8'b00010010;
		color_arr[9484] = 8'b00010010;
		color_arr[9485] = 8'b00010010;
		color_arr[9486] = 8'b00010010;
		color_arr[9487] = 8'b00010010;
		color_arr[9488] = 8'b00010010;
		color_arr[9489] = 8'b00010010;
		color_arr[9490] = 8'b00100000;
		color_arr[9491] = 8'b00100000;
		color_arr[9492] = 8'b00100000;
		color_arr[9493] = 8'b00000000;
		color_arr[9494] = 8'b00000000;
		color_arr[9495] = 8'b00100000;
		color_arr[9496] = 8'b00100000;
		color_arr[9497] = 8'b00100000;
		color_arr[9498] = 8'b00100000;
		color_arr[9499] = 8'b00100000;
		color_arr[9500] = 8'b00100000;
		color_arr[9501] = 8'b00100000;
		color_arr[9502] = 8'b00100000;
		color_arr[9503] = 8'b00100000;
		color_arr[9504] = 8'b00100000;
		color_arr[9505] = 8'b00100000;
		color_arr[9506] = 8'b00100000;
		color_arr[9507] = 8'b00100000;
		color_arr[9508] = 8'b00100000;
		color_arr[9509] = 8'b00100000;
		color_arr[9510] = 8'b00100000;
		color_arr[9511] = 8'b00100000;
		color_arr[9512] = 8'b00100000;
		color_arr[9513] = 8'b00100000;
		color_arr[9514] = 8'b00100000;
		color_arr[9515] = 8'b00100000;
		color_arr[9516] = 8'b00100000;
		color_arr[9517] = 8'b00100000;
		color_arr[9518] = 8'b00100000;
		color_arr[9519] = 8'b00100000;
		color_arr[9520] = 8'b00100000;
		color_arr[9521] = 8'b00100000;
		color_arr[9522] = 8'b00100000;
		color_arr[9523] = 8'b00100000;
		color_arr[9524] = 8'b00100000;
		color_arr[9525] = 8'b00100000;
		color_arr[9526] = 8'b00100000;
		color_arr[9527] = 8'b00100000;
		color_arr[9528] = 8'b00100000;
		color_arr[9529] = 8'b00100000;
		color_arr[9530] = 8'b00100000;
		color_arr[9531] = 8'b00100000;
		color_arr[9532] = 8'b00100000;
		color_arr[9533] = 8'b00100000;
		color_arr[9534] = 8'b00100000;
		color_arr[9535] = 8'b00100000;
		color_arr[9536] = 8'b00100000;
		color_arr[9537] = 8'b00100000;
		color_arr[9538] = 8'b00100000;
		color_arr[9539] = 8'b00100000;
		color_arr[9540] = 8'b00100000;
		color_arr[9541] = 8'b00100000;
		color_arr[9542] = 8'b00100000;
		color_arr[9543] = 8'b00100000;
		color_arr[9544] = 8'b00100000;
		color_arr[9545] = 8'b00100000;
		color_arr[9546] = 8'b00100000;
		color_arr[9547] = 8'b00100000;
		color_arr[9548] = 8'b00100000;
		color_arr[9549] = 8'b00100000;
		color_arr[9550] = 8'b00100000;
		color_arr[9551] = 8'b00100000;
		color_arr[9552] = 8'b00001000;
		color_arr[9553] = 8'b00001000;
		color_arr[9554] = 8'b00001000;
		color_arr[9555] = 8'b00001000;
		color_arr[9556] = 8'b00000000;
		color_arr[9557] = 8'b00000000;
		color_arr[9558] = 8'b00000000;
		color_arr[9559] = 8'b00001000;
		color_arr[9560] = 8'b00001000;
		color_arr[9561] = 8'b00001000;
		color_arr[9562] = 8'b00001000;
		color_arr[9563] = 8'b00001000;
		color_arr[9564] = 8'b00001000;
		color_arr[9565] = 8'b00001000;
		color_arr[9566] = 8'b00001000;
		color_arr[9567] = 8'b00001000;
		color_arr[9568] = 8'b00001000;
		color_arr[9569] = 8'b00001000;
		color_arr[9570] = 8'b00001000;
		color_arr[9571] = 8'b00001000;
		color_arr[9572] = 8'b00001000;
		color_arr[9573] = 8'b00001000;
		color_arr[9574] = 8'b00001000;
		color_arr[9575] = 8'b00001000;
		color_arr[9576] = 8'b00001000;
		color_arr[9577] = 8'b00001000;
		color_arr[9578] = 8'b00001000;
		color_arr[9579] = 8'b00001000;
		color_arr[9580] = 8'b00001000;
		color_arr[9581] = 8'b00001000;
		color_arr[9582] = 8'b00001000;
		color_arr[9583] = 8'b00001000;
		color_arr[9584] = 8'b00001000;
		color_arr[9585] = 8'b00001000;
		color_arr[9586] = 8'b00001000;
		color_arr[9587] = 8'b00001000;
		color_arr[9588] = 8'b00001000;
		color_arr[9589] = 8'b00000000;
		color_arr[9590] = 8'b00000000;
		color_arr[9591] = 8'b00000000;
		color_arr[9592] = 8'b00000000;
		color_arr[9593] = 8'b00001000;
		color_arr[9594] = 8'b00001000;
		color_arr[9595] = 8'b00001000;
		color_arr[9596] = 8'b00001000;
		color_arr[9597] = 8'b00010010;
		color_arr[9598] = 8'b00010010;
		color_arr[9599] = 8'b00010010;
		color_arr[9600] = 8'b00010010;
		color_arr[9601] = 8'b00010010;
		color_arr[9602] = 8'b00000000;
		color_arr[9603] = 8'b00000000;
		color_arr[9604] = 8'b00010010;
		color_arr[9605] = 8'b00010010;
		color_arr[9606] = 8'b00010010;
		color_arr[9607] = 8'b00010010;
		color_arr[9608] = 8'b00010010;
		color_arr[9609] = 8'b00010010;
		color_arr[9610] = 8'b00010010;
		color_arr[9611] = 8'b00010010;
		color_arr[9612] = 8'b00010010;
		color_arr[9613] = 8'b00010010;
		color_arr[9614] = 8'b00010010;
		color_arr[9615] = 8'b00010010;
		color_arr[9616] = 8'b00010010;
		color_arr[9617] = 8'b00010010;
		color_arr[9618] = 8'b00100000;
		color_arr[9619] = 8'b00100000;
		color_arr[9620] = 8'b00100000;
		color_arr[9621] = 8'b00000000;
		color_arr[9622] = 8'b00000000;
		color_arr[9623] = 8'b00100000;
		color_arr[9624] = 8'b00100000;
		color_arr[9625] = 8'b00100000;
		color_arr[9626] = 8'b00100000;
		color_arr[9627] = 8'b00100000;
		color_arr[9628] = 8'b00100000;
		color_arr[9629] = 8'b00100000;
		color_arr[9630] = 8'b00100000;
		color_arr[9631] = 8'b00100000;
		color_arr[9632] = 8'b00100000;
		color_arr[9633] = 8'b00100000;
		color_arr[9634] = 8'b00100000;
		color_arr[9635] = 8'b00100000;
		color_arr[9636] = 8'b00100000;
		color_arr[9637] = 8'b00100000;
		color_arr[9638] = 8'b00100000;
		color_arr[9639] = 8'b00100000;
		color_arr[9640] = 8'b00100000;
		color_arr[9641] = 8'b00100000;
		color_arr[9642] = 8'b00100000;
		color_arr[9643] = 8'b00100000;
		color_arr[9644] = 8'b00100000;
		color_arr[9645] = 8'b00100000;
		color_arr[9646] = 8'b00100000;
		color_arr[9647] = 8'b00100000;
		color_arr[9648] = 8'b00100000;
		color_arr[9649] = 8'b00100000;
		color_arr[9650] = 8'b00100000;
		color_arr[9651] = 8'b00100000;
		color_arr[9652] = 8'b00100000;
		color_arr[9653] = 8'b00100000;
		color_arr[9654] = 8'b00100000;
		color_arr[9655] = 8'b00100000;
		color_arr[9656] = 8'b00100000;
		color_arr[9657] = 8'b00100000;
		color_arr[9658] = 8'b00100000;
		color_arr[9659] = 8'b00100000;
		color_arr[9660] = 8'b00100000;
		color_arr[9661] = 8'b00100000;
		color_arr[9662] = 8'b00100000;
		color_arr[9663] = 8'b00100000;
		color_arr[9664] = 8'b00100000;
		color_arr[9665] = 8'b00100000;
		color_arr[9666] = 8'b00100000;
		color_arr[9667] = 8'b00100000;
		color_arr[9668] = 8'b00100000;
		color_arr[9669] = 8'b00100000;
		color_arr[9670] = 8'b00100000;
		color_arr[9671] = 8'b00100000;
		color_arr[9672] = 8'b00100000;
		color_arr[9673] = 8'b00100000;
		color_arr[9674] = 8'b00100000;
		color_arr[9675] = 8'b00100000;
		color_arr[9676] = 8'b00100000;
		color_arr[9677] = 8'b00100000;
		color_arr[9678] = 8'b00100000;
		color_arr[9679] = 8'b00100000;
		color_arr[9680] = 8'b00001000;
		color_arr[9681] = 8'b00001000;
		color_arr[9682] = 8'b00001000;
		color_arr[9683] = 8'b00001000;
		color_arr[9684] = 8'b00000000;
		color_arr[9685] = 8'b00000000;
		color_arr[9686] = 8'b00001000;
		color_arr[9687] = 8'b00001000;
		color_arr[9688] = 8'b00001000;
		color_arr[9689] = 8'b00001000;
		color_arr[9690] = 8'b00001000;
		color_arr[9691] = 8'b00001000;
		color_arr[9692] = 8'b00001000;
		color_arr[9693] = 8'b00001000;
		color_arr[9694] = 8'b00001000;
		color_arr[9695] = 8'b00001000;
		color_arr[9696] = 8'b00001000;
		color_arr[9697] = 8'b00001000;
		color_arr[9698] = 8'b00001000;
		color_arr[9699] = 8'b00001000;
		color_arr[9700] = 8'b00001000;
		color_arr[9701] = 8'b00001000;
		color_arr[9702] = 8'b00001000;
		color_arr[9703] = 8'b00001000;
		color_arr[9704] = 8'b00001000;
		color_arr[9705] = 8'b00001000;
		color_arr[9706] = 8'b00001000;
		color_arr[9707] = 8'b00001000;
		color_arr[9708] = 8'b00001000;
		color_arr[9709] = 8'b00001000;
		color_arr[9710] = 8'b00001000;
		color_arr[9711] = 8'b00001000;
		color_arr[9712] = 8'b00001000;
		color_arr[9713] = 8'b00001000;
		color_arr[9714] = 8'b00001000;
		color_arr[9715] = 8'b00001000;
		color_arr[9716] = 8'b00001000;
		color_arr[9717] = 8'b00000000;
		color_arr[9718] = 8'b00000000;
		color_arr[9719] = 8'b00000000;
		color_arr[9720] = 8'b00000000;
		color_arr[9721] = 8'b00001000;
		color_arr[9722] = 8'b00001000;
		color_arr[9723] = 8'b00001000;
		color_arr[9724] = 8'b00001000;
		color_arr[9725] = 8'b00010010;
		color_arr[9726] = 8'b00010010;
		color_arr[9727] = 8'b00010010;
		color_arr[9728] = 8'b00010010;
		color_arr[9729] = 8'b00010010;
		color_arr[9730] = 8'b00000000;
		color_arr[9731] = 8'b00000000;
		color_arr[9732] = 8'b00010010;
		color_arr[9733] = 8'b00010010;
		color_arr[9734] = 8'b00010010;
		color_arr[9735] = 8'b00010010;
		color_arr[9736] = 8'b00010010;
		color_arr[9737] = 8'b00010010;
		color_arr[9738] = 8'b00010010;
		color_arr[9739] = 8'b00010010;
		color_arr[9740] = 8'b00010010;
		color_arr[9741] = 8'b00010010;
		color_arr[9742] = 8'b00010010;
		color_arr[9743] = 8'b00010010;
		color_arr[9744] = 8'b00010010;
		color_arr[9745] = 8'b00010010;
		color_arr[9746] = 8'b00100000;
		color_arr[9747] = 8'b00100000;
		color_arr[9748] = 8'b00100000;
		color_arr[9749] = 8'b00000000;
		color_arr[9750] = 8'b00000000;
		color_arr[9751] = 8'b00100000;
		color_arr[9752] = 8'b00100000;
		color_arr[9753] = 8'b00100000;
		color_arr[9754] = 8'b00100000;
		color_arr[9755] = 8'b00100000;
		color_arr[9756] = 8'b00100000;
		color_arr[9757] = 8'b00100000;
		color_arr[9758] = 8'b00100000;
		color_arr[9759] = 8'b00100000;
		color_arr[9760] = 8'b00100000;
		color_arr[9761] = 8'b00100000;
		color_arr[9762] = 8'b00100000;
		color_arr[9763] = 8'b00100000;
		color_arr[9764] = 8'b00100000;
		color_arr[9765] = 8'b00100000;
		color_arr[9766] = 8'b00100000;
		color_arr[9767] = 8'b00100000;
		color_arr[9768] = 8'b00100000;
		color_arr[9769] = 8'b00100000;
		color_arr[9770] = 8'b00100000;
		color_arr[9771] = 8'b00100000;
		color_arr[9772] = 8'b00100000;
		color_arr[9773] = 8'b00100000;
		color_arr[9774] = 8'b00100000;
		color_arr[9775] = 8'b00100000;
		color_arr[9776] = 8'b00100000;
		color_arr[9777] = 8'b00100000;
		color_arr[9778] = 8'b00100000;
		color_arr[9779] = 8'b00100000;
		color_arr[9780] = 8'b00100000;
		color_arr[9781] = 8'b00100000;
		color_arr[9782] = 8'b00100000;
		color_arr[9783] = 8'b00100000;
		color_arr[9784] = 8'b00100000;
		color_arr[9785] = 8'b00100000;
		color_arr[9786] = 8'b00100000;
		color_arr[9787] = 8'b00100000;
		color_arr[9788] = 8'b00100000;
		color_arr[9789] = 8'b00100000;
		color_arr[9790] = 8'b00100000;
		color_arr[9791] = 8'b00100000;
		color_arr[9792] = 8'b00100000;
		color_arr[9793] = 8'b00100000;
		color_arr[9794] = 8'b00100000;
		color_arr[9795] = 8'b00100000;
		color_arr[9796] = 8'b00100000;
		color_arr[9797] = 8'b00100000;
		color_arr[9798] = 8'b00100000;
		color_arr[9799] = 8'b00100000;
		color_arr[9800] = 8'b00100000;
		color_arr[9801] = 8'b00100000;
		color_arr[9802] = 8'b00100000;
		color_arr[9803] = 8'b00100000;
		color_arr[9804] = 8'b00100000;
		color_arr[9805] = 8'b00100000;
		color_arr[9806] = 8'b00100000;
		color_arr[9807] = 8'b00100000;
		color_arr[9808] = 8'b00001000;
		color_arr[9809] = 8'b00001000;
		color_arr[9810] = 8'b00001000;
		color_arr[9811] = 8'b00000000;
		color_arr[9812] = 8'b00000000;
		color_arr[9813] = 8'b00000000;
		color_arr[9814] = 8'b00001000;
		color_arr[9815] = 8'b00001000;
		color_arr[9816] = 8'b00001000;
		color_arr[9817] = 8'b00001000;
		color_arr[9818] = 8'b00001000;
		color_arr[9819] = 8'b00001000;
		color_arr[9820] = 8'b00001000;
		color_arr[9821] = 8'b00001000;
		color_arr[9822] = 8'b00001000;
		color_arr[9823] = 8'b00001000;
		color_arr[9824] = 8'b00001000;
		color_arr[9825] = 8'b00001000;
		color_arr[9826] = 8'b00001000;
		color_arr[9827] = 8'b00001000;
		color_arr[9828] = 8'b00001000;
		color_arr[9829] = 8'b00001000;
		color_arr[9830] = 8'b00001000;
		color_arr[9831] = 8'b00001000;
		color_arr[9832] = 8'b00001000;
		color_arr[9833] = 8'b00001000;
		color_arr[9834] = 8'b00001000;
		color_arr[9835] = 8'b00001000;
		color_arr[9836] = 8'b00001000;
		color_arr[9837] = 8'b00001000;
		color_arr[9838] = 8'b00001000;
		color_arr[9839] = 8'b00001000;
		color_arr[9840] = 8'b00001000;
		color_arr[9841] = 8'b00001000;
		color_arr[9842] = 8'b00001000;
		color_arr[9843] = 8'b00001000;
		color_arr[9844] = 8'b00001000;
		color_arr[9845] = 8'b00000000;
		color_arr[9846] = 8'b00000000;
		color_arr[9847] = 8'b00000000;
		color_arr[9848] = 8'b00000000;
		color_arr[9849] = 8'b00001000;
		color_arr[9850] = 8'b00001000;
		color_arr[9851] = 8'b00001000;
		color_arr[9852] = 8'b00001000;
		color_arr[9853] = 8'b00010010;
		color_arr[9854] = 8'b00010010;
		color_arr[9855] = 8'b00010010;
		color_arr[9856] = 8'b00010010;
		color_arr[9857] = 8'b00010010;
		color_arr[9858] = 8'b00000000;
		color_arr[9859] = 8'b00000000;
		color_arr[9860] = 8'b00010010;
		color_arr[9861] = 8'b00010010;
		color_arr[9862] = 8'b00010010;
		color_arr[9863] = 8'b00010010;
		color_arr[9864] = 8'b00010010;
		color_arr[9865] = 8'b00010010;
		color_arr[9866] = 8'b00010010;
		color_arr[9867] = 8'b00010010;
		color_arr[9868] = 8'b00010010;
		color_arr[9869] = 8'b00010010;
		color_arr[9870] = 8'b00010010;
		color_arr[9871] = 8'b00010010;
		color_arr[9872] = 8'b00010010;
		color_arr[9873] = 8'b00010010;
		color_arr[9874] = 8'b00100000;
		color_arr[9875] = 8'b00100000;
		color_arr[9876] = 8'b00100000;
		color_arr[9877] = 8'b00000000;
		color_arr[9878] = 8'b00000000;
		color_arr[9879] = 8'b00100000;
		color_arr[9880] = 8'b00100000;
		color_arr[9881] = 8'b00100000;
		color_arr[9882] = 8'b00100000;
		color_arr[9883] = 8'b00100000;
		color_arr[9884] = 8'b00100000;
		color_arr[9885] = 8'b00100000;
		color_arr[9886] = 8'b00100000;
		color_arr[9887] = 8'b00100000;
		color_arr[9888] = 8'b00100000;
		color_arr[9889] = 8'b00100000;
		color_arr[9890] = 8'b00100000;
		color_arr[9891] = 8'b00100000;
		color_arr[9892] = 8'b00100000;
		color_arr[9893] = 8'b00100000;
		color_arr[9894] = 8'b00100000;
		color_arr[9895] = 8'b00100000;
		color_arr[9896] = 8'b00100000;
		color_arr[9897] = 8'b00100000;
		color_arr[9898] = 8'b00100000;
		color_arr[9899] = 8'b00100000;
		color_arr[9900] = 8'b00100000;
		color_arr[9901] = 8'b00100000;
		color_arr[9902] = 8'b00100000;
		color_arr[9903] = 8'b00100000;
		color_arr[9904] = 8'b00100000;
		color_arr[9905] = 8'b00100000;
		color_arr[9906] = 8'b00100000;
		color_arr[9907] = 8'b00100000;
		color_arr[9908] = 8'b00100000;
		color_arr[9909] = 8'b00100000;
		color_arr[9910] = 8'b00100000;
		color_arr[9911] = 8'b00100000;
		color_arr[9912] = 8'b00100000;
		color_arr[9913] = 8'b00100000;
		color_arr[9914] = 8'b00100000;
		color_arr[9915] = 8'b00100000;
		color_arr[9916] = 8'b00100000;
		color_arr[9917] = 8'b00100000;
		color_arr[9918] = 8'b00100000;
		color_arr[9919] = 8'b00100000;
		color_arr[9920] = 8'b00100000;
		color_arr[9921] = 8'b00100000;
		color_arr[9922] = 8'b00100000;
		color_arr[9923] = 8'b00100000;
		color_arr[9924] = 8'b00100000;
		color_arr[9925] = 8'b00100000;
		color_arr[9926] = 8'b00100000;
		color_arr[9927] = 8'b00100000;
		color_arr[9928] = 8'b00100000;
		color_arr[9929] = 8'b00100000;
		color_arr[9930] = 8'b00100000;
		color_arr[9931] = 8'b00100000;
		color_arr[9932] = 8'b00100000;
		color_arr[9933] = 8'b00100000;
		color_arr[9934] = 8'b00100000;
		color_arr[9935] = 8'b00100000;
		color_arr[9936] = 8'b00001000;
		color_arr[9937] = 8'b00001000;
		color_arr[9938] = 8'b00000000;
		color_arr[9939] = 8'b00000000;
		color_arr[9940] = 8'b00000000;
		color_arr[9941] = 8'b00001000;
		color_arr[9942] = 8'b00001000;
		color_arr[9943] = 8'b00001000;
		color_arr[9944] = 8'b00001000;
		color_arr[9945] = 8'b00001000;
		color_arr[9946] = 8'b00001000;
		color_arr[9947] = 8'b00001000;
		color_arr[9948] = 8'b00001000;
		color_arr[9949] = 8'b00001000;
		color_arr[9950] = 8'b00001000;
		color_arr[9951] = 8'b00001000;
		color_arr[9952] = 8'b00001000;
		color_arr[9953] = 8'b00001000;
		color_arr[9954] = 8'b00001000;
		color_arr[9955] = 8'b00001000;
		color_arr[9956] = 8'b00001000;
		color_arr[9957] = 8'b00001000;
		color_arr[9958] = 8'b00001000;
		color_arr[9959] = 8'b00001000;
		color_arr[9960] = 8'b00001000;
		color_arr[9961] = 8'b00001000;
		color_arr[9962] = 8'b00001000;
		color_arr[9963] = 8'b00001000;
		color_arr[9964] = 8'b00001000;
		color_arr[9965] = 8'b00001000;
		color_arr[9966] = 8'b00001000;
		color_arr[9967] = 8'b00001000;
		color_arr[9968] = 8'b00001000;
		color_arr[9969] = 8'b00001000;
		color_arr[9970] = 8'b00001000;
		color_arr[9971] = 8'b00001000;
		color_arr[9972] = 8'b00001000;
		color_arr[9973] = 8'b00000000;
		color_arr[9974] = 8'b00000000;
		color_arr[9975] = 8'b00000000;
		color_arr[9976] = 8'b00000000;
		color_arr[9977] = 8'b00001000;
		color_arr[9978] = 8'b00001000;
		color_arr[9979] = 8'b00001000;
		color_arr[9980] = 8'b00001000;
		color_arr[9981] = 8'b00010010;
		color_arr[9982] = 8'b00010010;
		color_arr[9983] = 8'b00010010;
		color_arr[9984] = 8'b00010010;
		color_arr[9985] = 8'b00010010;
		color_arr[9986] = 8'b00000000;
		color_arr[9987] = 8'b00000000;
		color_arr[9988] = 8'b00010010;
		color_arr[9989] = 8'b00010010;
		color_arr[9990] = 8'b00010010;
		color_arr[9991] = 8'b00010010;
		color_arr[9992] = 8'b00010010;
		color_arr[9993] = 8'b00010010;
		color_arr[9994] = 8'b00010010;
		color_arr[9995] = 8'b00010010;
		color_arr[9996] = 8'b00010010;
		color_arr[9997] = 8'b00010010;
		color_arr[9998] = 8'b00010010;
		color_arr[9999] = 8'b00010010;
		color_arr[10000] = 8'b00010010;
		color_arr[10001] = 8'b00010010;
		color_arr[10002] = 8'b00100000;
		color_arr[10003] = 8'b00100000;
		color_arr[10004] = 8'b00100000;
		color_arr[10005] = 8'b00000000;
		color_arr[10006] = 8'b00000000;
		color_arr[10007] = 8'b00100000;
		color_arr[10008] = 8'b00100000;
		color_arr[10009] = 8'b00100000;
		color_arr[10010] = 8'b00100000;
		color_arr[10011] = 8'b00100000;
		color_arr[10012] = 8'b00100000;
		color_arr[10013] = 8'b00100000;
		color_arr[10014] = 8'b00100000;
		color_arr[10015] = 8'b00100000;
		color_arr[10016] = 8'b00100000;
		color_arr[10017] = 8'b00100000;
		color_arr[10018] = 8'b00100000;
		color_arr[10019] = 8'b00100000;
		color_arr[10020] = 8'b00100000;
		color_arr[10021] = 8'b00100000;
		color_arr[10022] = 8'b00100000;
		color_arr[10023] = 8'b00100000;
		color_arr[10024] = 8'b00100000;
		color_arr[10025] = 8'b00100000;
		color_arr[10026] = 8'b00100000;
		color_arr[10027] = 8'b00100000;
		color_arr[10028] = 8'b00100000;
		color_arr[10029] = 8'b00100000;
		color_arr[10030] = 8'b00100000;
		color_arr[10031] = 8'b00100000;
		color_arr[10032] = 8'b00100000;
		color_arr[10033] = 8'b00100000;
		color_arr[10034] = 8'b00100000;
		color_arr[10035] = 8'b00100000;
		color_arr[10036] = 8'b00100000;
		color_arr[10037] = 8'b00100000;
		color_arr[10038] = 8'b00100000;
		color_arr[10039] = 8'b00100000;
		color_arr[10040] = 8'b00100000;
		color_arr[10041] = 8'b00100000;
		color_arr[10042] = 8'b00100000;
		color_arr[10043] = 8'b00100000;
		color_arr[10044] = 8'b00100000;
		color_arr[10045] = 8'b00100000;
		color_arr[10046] = 8'b00100000;
		color_arr[10047] = 8'b00100000;
		color_arr[10048] = 8'b00100000;
		color_arr[10049] = 8'b00100000;
		color_arr[10050] = 8'b00100000;
		color_arr[10051] = 8'b00100000;
		color_arr[10052] = 8'b00100000;
		color_arr[10053] = 8'b00100000;
		color_arr[10054] = 8'b00100000;
		color_arr[10055] = 8'b00100000;
		color_arr[10056] = 8'b00100000;
		color_arr[10057] = 8'b00100000;
		color_arr[10058] = 8'b00100000;
		color_arr[10059] = 8'b00100000;
		color_arr[10060] = 8'b00100000;
		color_arr[10061] = 8'b00100000;
		color_arr[10062] = 8'b00100000;
		color_arr[10063] = 8'b00100000;
		color_arr[10064] = 8'b00001000;
		color_arr[10065] = 8'b00000000;
		color_arr[10066] = 8'b00000000;
		color_arr[10067] = 8'b00000000;
		color_arr[10068] = 8'b00001000;
		color_arr[10069] = 8'b00001000;
		color_arr[10070] = 8'b00001000;
		color_arr[10071] = 8'b00001000;
		color_arr[10072] = 8'b00001000;
		color_arr[10073] = 8'b00001000;
		color_arr[10074] = 8'b00001000;
		color_arr[10075] = 8'b00001000;
		color_arr[10076] = 8'b00001000;
		color_arr[10077] = 8'b00001000;
		color_arr[10078] = 8'b00001000;
		color_arr[10079] = 8'b00001000;
		color_arr[10080] = 8'b00001000;
		color_arr[10081] = 8'b00001000;
		color_arr[10082] = 8'b00001000;
		color_arr[10083] = 8'b00001000;
		color_arr[10084] = 8'b00001000;
		color_arr[10085] = 8'b00001000;
		color_arr[10086] = 8'b00001000;
		color_arr[10087] = 8'b00001000;
		color_arr[10088] = 8'b00001000;
		color_arr[10089] = 8'b00001000;
		color_arr[10090] = 8'b00001000;
		color_arr[10091] = 8'b00001000;
		color_arr[10092] = 8'b00001000;
		color_arr[10093] = 8'b00001000;
		color_arr[10094] = 8'b00001000;
		color_arr[10095] = 8'b00001000;
		color_arr[10096] = 8'b00001000;
		color_arr[10097] = 8'b00001000;
		color_arr[10098] = 8'b00001000;
		color_arr[10099] = 8'b00001000;
		color_arr[10100] = 8'b00001000;
		color_arr[10101] = 8'b00000000;
		color_arr[10102] = 8'b00000000;
		color_arr[10103] = 8'b00000000;
		color_arr[10104] = 8'b00000000;
		color_arr[10105] = 8'b00001000;
		color_arr[10106] = 8'b00001000;
		color_arr[10107] = 8'b00001000;
		color_arr[10108] = 8'b00001000;
		color_arr[10109] = 8'b00010010;
		color_arr[10110] = 8'b00010010;
		color_arr[10111] = 8'b00010010;
		color_arr[10112] = 8'b00010010;
		color_arr[10113] = 8'b00010010;
		color_arr[10114] = 8'b00000000;
		color_arr[10115] = 8'b00000000;
		color_arr[10116] = 8'b00010010;
		color_arr[10117] = 8'b00010010;
		color_arr[10118] = 8'b00010010;
		color_arr[10119] = 8'b00010010;
		color_arr[10120] = 8'b00010010;
		color_arr[10121] = 8'b00010010;
		color_arr[10122] = 8'b00010010;
		color_arr[10123] = 8'b00010010;
		color_arr[10124] = 8'b00010010;
		color_arr[10125] = 8'b00010010;
		color_arr[10126] = 8'b00010010;
		color_arr[10127] = 8'b00010010;
		color_arr[10128] = 8'b00010010;
		color_arr[10129] = 8'b00010010;
		color_arr[10130] = 8'b00100000;
		color_arr[10131] = 8'b00100000;
		color_arr[10132] = 8'b00100000;
		color_arr[10133] = 8'b00000000;
		color_arr[10134] = 8'b00000000;
		color_arr[10135] = 8'b00000000;
		color_arr[10136] = 8'b00100000;
		color_arr[10137] = 8'b00100000;
		color_arr[10138] = 8'b00100000;
		color_arr[10139] = 8'b00100000;
		color_arr[10140] = 8'b00100000;
		color_arr[10141] = 8'b00100000;
		color_arr[10142] = 8'b00100000;
		color_arr[10143] = 8'b00100000;
		color_arr[10144] = 8'b00100000;
		color_arr[10145] = 8'b00100000;
		color_arr[10146] = 8'b00100000;
		color_arr[10147] = 8'b00100000;
		color_arr[10148] = 8'b00100000;
		color_arr[10149] = 8'b00100000;
		color_arr[10150] = 8'b00100000;
		color_arr[10151] = 8'b00100000;
		color_arr[10152] = 8'b00100000;
		color_arr[10153] = 8'b00100000;
		color_arr[10154] = 8'b00100000;
		color_arr[10155] = 8'b00100000;
		color_arr[10156] = 8'b00100000;
		color_arr[10157] = 8'b00100000;
		color_arr[10158] = 8'b00100000;
		color_arr[10159] = 8'b00100000;
		color_arr[10160] = 8'b00100000;
		color_arr[10161] = 8'b00100000;
		color_arr[10162] = 8'b00100000;
		color_arr[10163] = 8'b00100000;
		color_arr[10164] = 8'b00100000;
		color_arr[10165] = 8'b00100000;
		color_arr[10166] = 8'b00100000;
		color_arr[10167] = 8'b00100000;
		color_arr[10168] = 8'b00100000;
		color_arr[10169] = 8'b00100000;
		color_arr[10170] = 8'b00100000;
		color_arr[10171] = 8'b00100000;
		color_arr[10172] = 8'b00100000;
		color_arr[10173] = 8'b00100000;
		color_arr[10174] = 8'b00100000;
		color_arr[10175] = 8'b00100000;
		color_arr[10176] = 8'b00100000;
		color_arr[10177] = 8'b00100000;
		color_arr[10178] = 8'b00100000;
		color_arr[10179] = 8'b00100000;
		color_arr[10180] = 8'b00100000;
		color_arr[10181] = 8'b00100000;
		color_arr[10182] = 8'b00100000;
		color_arr[10183] = 8'b00100000;
		color_arr[10184] = 8'b00100000;
		color_arr[10185] = 8'b00100000;
		color_arr[10186] = 8'b00100000;
		color_arr[10187] = 8'b00100000;
		color_arr[10188] = 8'b00100000;
		color_arr[10189] = 8'b00100000;
		color_arr[10190] = 8'b00100000;
		color_arr[10191] = 8'b00100000;
		color_arr[10192] = 8'b00000000;
		color_arr[10193] = 8'b00000000;
		color_arr[10194] = 8'b00000000;
		color_arr[10195] = 8'b00001000;
		color_arr[10196] = 8'b00001000;
		color_arr[10197] = 8'b00001000;
		color_arr[10198] = 8'b00001000;
		color_arr[10199] = 8'b00001000;
		color_arr[10200] = 8'b00001000;
		color_arr[10201] = 8'b00001000;
		color_arr[10202] = 8'b00001000;
		color_arr[10203] = 8'b00001000;
		color_arr[10204] = 8'b00001000;
		color_arr[10205] = 8'b00001000;
		color_arr[10206] = 8'b00001000;
		color_arr[10207] = 8'b00001000;
		color_arr[10208] = 8'b00001000;
		color_arr[10209] = 8'b00001000;
		color_arr[10210] = 8'b00001000;
		color_arr[10211] = 8'b00001000;
		color_arr[10212] = 8'b00001000;
		color_arr[10213] = 8'b00001000;
		color_arr[10214] = 8'b00001000;
		color_arr[10215] = 8'b00001000;
		color_arr[10216] = 8'b00001000;
		color_arr[10217] = 8'b00001000;
		color_arr[10218] = 8'b00001000;
		color_arr[10219] = 8'b00001000;
		color_arr[10220] = 8'b00001000;
		color_arr[10221] = 8'b00001000;
		color_arr[10222] = 8'b00001000;
		color_arr[10223] = 8'b00001000;
		color_arr[10224] = 8'b00001000;
		color_arr[10225] = 8'b00001000;
		color_arr[10226] = 8'b00001000;
		color_arr[10227] = 8'b00001000;
		color_arr[10228] = 8'b00001000;
		color_arr[10229] = 8'b00000000;
		color_arr[10230] = 8'b00000000;
		color_arr[10231] = 8'b00000000;
		color_arr[10232] = 8'b00000000;
		color_arr[10233] = 8'b00001000;
		color_arr[10234] = 8'b00001000;
		color_arr[10235] = 8'b00001000;
		color_arr[10236] = 8'b00001000;
		color_arr[10237] = 8'b00010010;
		color_arr[10238] = 8'b00010010;
		color_arr[10239] = 8'b00010010;
		color_arr[10240] = 8'b00010010;
		color_arr[10241] = 8'b00010010;
		color_arr[10242] = 8'b00000000;
		color_arr[10243] = 8'b00000000;
		color_arr[10244] = 8'b00010010;
		color_arr[10245] = 8'b00010010;
		color_arr[10246] = 8'b00010010;
		color_arr[10247] = 8'b00010010;
		color_arr[10248] = 8'b00010010;
		color_arr[10249] = 8'b00010010;
		color_arr[10250] = 8'b00010010;
		color_arr[10251] = 8'b00010010;
		color_arr[10252] = 8'b00010010;
		color_arr[10253] = 8'b00010010;
		color_arr[10254] = 8'b00010010;
		color_arr[10255] = 8'b00010010;
		color_arr[10256] = 8'b00010010;
		color_arr[10257] = 8'b00010010;
		color_arr[10258] = 8'b00100000;
		color_arr[10259] = 8'b00100000;
		color_arr[10260] = 8'b00100000;
		color_arr[10261] = 8'b00100000;
		color_arr[10262] = 8'b00000000;
		color_arr[10263] = 8'b00000000;
		color_arr[10264] = 8'b00100000;
		color_arr[10265] = 8'b00100000;
		color_arr[10266] = 8'b00100000;
		color_arr[10267] = 8'b00100000;
		color_arr[10268] = 8'b00100000;
		color_arr[10269] = 8'b00100000;
		color_arr[10270] = 8'b00100000;
		color_arr[10271] = 8'b00100000;
		color_arr[10272] = 8'b00100000;
		color_arr[10273] = 8'b00100000;
		color_arr[10274] = 8'b00100000;
		color_arr[10275] = 8'b00100000;
		color_arr[10276] = 8'b00100000;
		color_arr[10277] = 8'b00100000;
		color_arr[10278] = 8'b00100000;
		color_arr[10279] = 8'b00100000;
		color_arr[10280] = 8'b00100000;
		color_arr[10281] = 8'b00100000;
		color_arr[10282] = 8'b00100000;
		color_arr[10283] = 8'b00100000;
		color_arr[10284] = 8'b00100000;
		color_arr[10285] = 8'b00100000;
		color_arr[10286] = 8'b00100000;
		color_arr[10287] = 8'b00100000;
		color_arr[10288] = 8'b00100000;
		color_arr[10289] = 8'b00100000;
		color_arr[10290] = 8'b00100000;
		color_arr[10291] = 8'b00100000;
		color_arr[10292] = 8'b00100000;
		color_arr[10293] = 8'b00100000;
		color_arr[10294] = 8'b00100000;
		color_arr[10295] = 8'b00100000;
		color_arr[10296] = 8'b00100000;
		color_arr[10297] = 8'b00100000;
		color_arr[10298] = 8'b00100000;
		color_arr[10299] = 8'b00100000;
		color_arr[10300] = 8'b00100000;
		color_arr[10301] = 8'b00100000;
		color_arr[10302] = 8'b00100000;
		color_arr[10303] = 8'b00100000;
		color_arr[10304] = 8'b00100000;
		color_arr[10305] = 8'b00100000;
		color_arr[10306] = 8'b00100000;
		color_arr[10307] = 8'b00100000;
		color_arr[10308] = 8'b00100000;
		color_arr[10309] = 8'b00100000;
		color_arr[10310] = 8'b00100000;
		color_arr[10311] = 8'b00100000;
		color_arr[10312] = 8'b00100000;
		color_arr[10313] = 8'b00100000;
		color_arr[10314] = 8'b00100000;
		color_arr[10315] = 8'b00100000;
		color_arr[10316] = 8'b00100000;
		color_arr[10317] = 8'b00100000;
		color_arr[10318] = 8'b00100000;
		color_arr[10319] = 8'b00000000;
		color_arr[10320] = 8'b00000000;
		color_arr[10321] = 8'b00000000;
		color_arr[10322] = 8'b00001000;
		color_arr[10323] = 8'b00001000;
		color_arr[10324] = 8'b00001000;
		color_arr[10325] = 8'b00001000;
		color_arr[10326] = 8'b00001000;
		color_arr[10327] = 8'b00001000;
		color_arr[10328] = 8'b00001000;
		color_arr[10329] = 8'b00001000;
		color_arr[10330] = 8'b00001000;
		color_arr[10331] = 8'b00001000;
		color_arr[10332] = 8'b00001000;
		color_arr[10333] = 8'b00001000;
		color_arr[10334] = 8'b00001000;
		color_arr[10335] = 8'b00001000;
		color_arr[10336] = 8'b00001000;
		color_arr[10337] = 8'b00001000;
		color_arr[10338] = 8'b00001000;
		color_arr[10339] = 8'b00001000;
		color_arr[10340] = 8'b00001000;
		color_arr[10341] = 8'b00001000;
		color_arr[10342] = 8'b00001000;
		color_arr[10343] = 8'b00001000;
		color_arr[10344] = 8'b00001000;
		color_arr[10345] = 8'b00001000;
		color_arr[10346] = 8'b00001000;
		color_arr[10347] = 8'b00001000;
		color_arr[10348] = 8'b00001000;
		color_arr[10349] = 8'b00001000;
		color_arr[10350] = 8'b00001000;
		color_arr[10351] = 8'b00001000;
		color_arr[10352] = 8'b00001000;
		color_arr[10353] = 8'b00001000;
		color_arr[10354] = 8'b00001000;
		color_arr[10355] = 8'b00001000;
		color_arr[10356] = 8'b00001000;
		color_arr[10357] = 8'b00000000;
		color_arr[10358] = 8'b00000000;
		color_arr[10359] = 8'b00000000;
		color_arr[10360] = 8'b00000000;
		color_arr[10361] = 8'b00001000;
		color_arr[10362] = 8'b00001000;
		color_arr[10363] = 8'b00001000;
		color_arr[10364] = 8'b00001000;
		color_arr[10365] = 8'b00010010;
		color_arr[10366] = 8'b00010010;
		color_arr[10367] = 8'b00010010;
		color_arr[10368] = 8'b00010010;
		color_arr[10369] = 8'b00010010;
		color_arr[10370] = 8'b00000000;
		color_arr[10371] = 8'b00000000;
		color_arr[10372] = 8'b00010010;
		color_arr[10373] = 8'b00010010;
		color_arr[10374] = 8'b00010010;
		color_arr[10375] = 8'b00010010;
		color_arr[10376] = 8'b00010010;
		color_arr[10377] = 8'b00010010;
		color_arr[10378] = 8'b00010010;
		color_arr[10379] = 8'b00010010;
		color_arr[10380] = 8'b00010010;
		color_arr[10381] = 8'b00010010;
		color_arr[10382] = 8'b00010010;
		color_arr[10383] = 8'b00010010;
		color_arr[10384] = 8'b00010010;
		color_arr[10385] = 8'b00010010;
		color_arr[10386] = 8'b00100000;
		color_arr[10387] = 8'b00100000;
		color_arr[10388] = 8'b00100000;
		color_arr[10389] = 8'b00100000;
		color_arr[10390] = 8'b00000000;
		color_arr[10391] = 8'b00000000;
		color_arr[10392] = 8'b00100000;
		color_arr[10393] = 8'b00100000;
		color_arr[10394] = 8'b00100000;
		color_arr[10395] = 8'b00100000;
		color_arr[10396] = 8'b00100000;
		color_arr[10397] = 8'b00100000;
		color_arr[10398] = 8'b00100000;
		color_arr[10399] = 8'b00100000;
		color_arr[10400] = 8'b00100000;
		color_arr[10401] = 8'b00100000;
		color_arr[10402] = 8'b00100000;
		color_arr[10403] = 8'b00100000;
		color_arr[10404] = 8'b00100000;
		color_arr[10405] = 8'b00100000;
		color_arr[10406] = 8'b00100000;
		color_arr[10407] = 8'b00100000;
		color_arr[10408] = 8'b00100000;
		color_arr[10409] = 8'b00100000;
		color_arr[10410] = 8'b00100000;
		color_arr[10411] = 8'b00100000;
		color_arr[10412] = 8'b00100000;
		color_arr[10413] = 8'b00100000;
		color_arr[10414] = 8'b00100000;
		color_arr[10415] = 8'b00100000;
		color_arr[10416] = 8'b00100000;
		color_arr[10417] = 8'b00100000;
		color_arr[10418] = 8'b00100000;
		color_arr[10419] = 8'b00100000;
		color_arr[10420] = 8'b00100000;
		color_arr[10421] = 8'b00100000;
		color_arr[10422] = 8'b00100000;
		color_arr[10423] = 8'b00100000;
		color_arr[10424] = 8'b00100000;
		color_arr[10425] = 8'b00100000;
		color_arr[10426] = 8'b00100000;
		color_arr[10427] = 8'b00100000;
		color_arr[10428] = 8'b00100000;
		color_arr[10429] = 8'b00100000;
		color_arr[10430] = 8'b00100000;
		color_arr[10431] = 8'b00100000;
		color_arr[10432] = 8'b00100000;
		color_arr[10433] = 8'b00100000;
		color_arr[10434] = 8'b00100000;
		color_arr[10435] = 8'b00100000;
		color_arr[10436] = 8'b00100000;
		color_arr[10437] = 8'b00100000;
		color_arr[10438] = 8'b00100000;
		color_arr[10439] = 8'b00100000;
		color_arr[10440] = 8'b00100000;
		color_arr[10441] = 8'b00100000;
		color_arr[10442] = 8'b00100000;
		color_arr[10443] = 8'b00100000;
		color_arr[10444] = 8'b00100000;
		color_arr[10445] = 8'b00100000;
		color_arr[10446] = 8'b00100000;
		color_arr[10447] = 8'b00000000;
		color_arr[10448] = 8'b00000000;
		color_arr[10449] = 8'b00001000;
		color_arr[10450] = 8'b00001000;
		color_arr[10451] = 8'b00001000;
		color_arr[10452] = 8'b00001000;
		color_arr[10453] = 8'b00001000;
		color_arr[10454] = 8'b00001000;
		color_arr[10455] = 8'b00001000;
		color_arr[10456] = 8'b00001000;
		color_arr[10457] = 8'b00001000;
		color_arr[10458] = 8'b00001000;
		color_arr[10459] = 8'b00001000;
		color_arr[10460] = 8'b00001000;
		color_arr[10461] = 8'b00001000;
		color_arr[10462] = 8'b00001000;
		color_arr[10463] = 8'b00001000;
		color_arr[10464] = 8'b00001000;
		color_arr[10465] = 8'b00001000;
		color_arr[10466] = 8'b00001000;
		color_arr[10467] = 8'b00001000;
		color_arr[10468] = 8'b00001000;
		color_arr[10469] = 8'b00001000;
		color_arr[10470] = 8'b00001000;
		color_arr[10471] = 8'b00001000;
		color_arr[10472] = 8'b00001000;
		color_arr[10473] = 8'b00001000;
		color_arr[10474] = 8'b00001000;
		color_arr[10475] = 8'b00001000;
		color_arr[10476] = 8'b00001000;
		color_arr[10477] = 8'b00001000;
		color_arr[10478] = 8'b00001000;
		color_arr[10479] = 8'b00001000;
		color_arr[10480] = 8'b00001000;
		color_arr[10481] = 8'b00001000;
		color_arr[10482] = 8'b00001000;
		color_arr[10483] = 8'b00001000;
		color_arr[10484] = 8'b00001000;
		color_arr[10485] = 8'b00000000;
		color_arr[10486] = 8'b00000000;
		color_arr[10487] = 8'b00000000;
		color_arr[10488] = 8'b00000000;
		color_arr[10489] = 8'b00001000;
		color_arr[10490] = 8'b00001000;
		color_arr[10491] = 8'b00001000;
		color_arr[10492] = 8'b00001000;
		color_arr[10493] = 8'b00010010;
		color_arr[10494] = 8'b00010010;
		color_arr[10495] = 8'b00010010;
		color_arr[10496] = 8'b00010010;
		color_arr[10497] = 8'b00000000;
		color_arr[10498] = 8'b00000000;
		color_arr[10499] = 8'b00000000;
		color_arr[10500] = 8'b00010010;
		color_arr[10501] = 8'b00010010;
		color_arr[10502] = 8'b00010010;
		color_arr[10503] = 8'b00010010;
		color_arr[10504] = 8'b00010010;
		color_arr[10505] = 8'b00010010;
		color_arr[10506] = 8'b00010010;
		color_arr[10507] = 8'b00010010;
		color_arr[10508] = 8'b00010010;
		color_arr[10509] = 8'b00010010;
		color_arr[10510] = 8'b00010010;
		color_arr[10511] = 8'b00010010;
		color_arr[10512] = 8'b00010010;
		color_arr[10513] = 8'b00010010;
		color_arr[10514] = 8'b00100000;
		color_arr[10515] = 8'b00100000;
		color_arr[10516] = 8'b00100000;
		color_arr[10517] = 8'b00100000;
		color_arr[10518] = 8'b00000000;
		color_arr[10519] = 8'b00000000;
		color_arr[10520] = 8'b00100000;
		color_arr[10521] = 8'b00100000;
		color_arr[10522] = 8'b00100000;
		color_arr[10523] = 8'b00100000;
		color_arr[10524] = 8'b00100000;
		color_arr[10525] = 8'b00100000;
		color_arr[10526] = 8'b00100000;
		color_arr[10527] = 8'b00100000;
		color_arr[10528] = 8'b00100000;
		color_arr[10529] = 8'b00100000;
		color_arr[10530] = 8'b00100000;
		color_arr[10531] = 8'b00100000;
		color_arr[10532] = 8'b00100000;
		color_arr[10533] = 8'b00100000;
		color_arr[10534] = 8'b00100000;
		color_arr[10535] = 8'b00100000;
		color_arr[10536] = 8'b00100000;
		color_arr[10537] = 8'b00100000;
		color_arr[10538] = 8'b00100000;
		color_arr[10539] = 8'b00100000;
		color_arr[10540] = 8'b00100000;
		color_arr[10541] = 8'b00100000;
		color_arr[10542] = 8'b00100000;
		color_arr[10543] = 8'b00100000;
		color_arr[10544] = 8'b00100000;
		color_arr[10545] = 8'b00100000;
		color_arr[10546] = 8'b00100000;
		color_arr[10547] = 8'b00100000;
		color_arr[10548] = 8'b00100000;
		color_arr[10549] = 8'b00100000;
		color_arr[10550] = 8'b00100000;
		color_arr[10551] = 8'b00100000;
		color_arr[10552] = 8'b00100000;
		color_arr[10553] = 8'b00100000;
		color_arr[10554] = 8'b00100000;
		color_arr[10555] = 8'b00100000;
		color_arr[10556] = 8'b00100000;
		color_arr[10557] = 8'b00100000;
		color_arr[10558] = 8'b00100000;
		color_arr[10559] = 8'b00100000;
		color_arr[10560] = 8'b00100000;
		color_arr[10561] = 8'b00100000;
		color_arr[10562] = 8'b00100000;
		color_arr[10563] = 8'b00100000;
		color_arr[10564] = 8'b00100000;
		color_arr[10565] = 8'b00100000;
		color_arr[10566] = 8'b00100000;
		color_arr[10567] = 8'b00100000;
		color_arr[10568] = 8'b00100000;
		color_arr[10569] = 8'b00100000;
		color_arr[10570] = 8'b00100000;
		color_arr[10571] = 8'b00100000;
		color_arr[10572] = 8'b00100000;
		color_arr[10573] = 8'b00100000;
		color_arr[10574] = 8'b00000000;
		color_arr[10575] = 8'b00000000;
		color_arr[10576] = 8'b00000000;
		color_arr[10577] = 8'b00001000;
		color_arr[10578] = 8'b00001000;
		color_arr[10579] = 8'b00001000;
		color_arr[10580] = 8'b00001000;
		color_arr[10581] = 8'b00001000;
		color_arr[10582] = 8'b00001000;
		color_arr[10583] = 8'b00001000;
		color_arr[10584] = 8'b00001000;
		color_arr[10585] = 8'b00001000;
		color_arr[10586] = 8'b00001000;
		color_arr[10587] = 8'b00001000;
		color_arr[10588] = 8'b00001000;
		color_arr[10589] = 8'b00001000;
		color_arr[10590] = 8'b00001000;
		color_arr[10591] = 8'b00001000;
		color_arr[10592] = 8'b00001000;
		color_arr[10593] = 8'b00001000;
		color_arr[10594] = 8'b00001000;
		color_arr[10595] = 8'b00001000;
		color_arr[10596] = 8'b00001000;
		color_arr[10597] = 8'b00001000;
		color_arr[10598] = 8'b00001000;
		color_arr[10599] = 8'b00001000;
		color_arr[10600] = 8'b00001000;
		color_arr[10601] = 8'b00001000;
		color_arr[10602] = 8'b00001000;
		color_arr[10603] = 8'b00001000;
		color_arr[10604] = 8'b00001000;
		color_arr[10605] = 8'b00001000;
		color_arr[10606] = 8'b00001000;
		color_arr[10607] = 8'b00001000;
		color_arr[10608] = 8'b00001000;
		color_arr[10609] = 8'b00001000;
		color_arr[10610] = 8'b00001000;
		color_arr[10611] = 8'b00001000;
		color_arr[10612] = 8'b00001000;
		color_arr[10613] = 8'b00000000;
		color_arr[10614] = 8'b00000000;
		color_arr[10615] = 8'b00000000;
		color_arr[10616] = 8'b00000000;
		color_arr[10617] = 8'b00001000;
		color_arr[10618] = 8'b00001000;
		color_arr[10619] = 8'b00001000;
		color_arr[10620] = 8'b00001000;
		color_arr[10621] = 8'b00010010;
		color_arr[10622] = 8'b00010010;
		color_arr[10623] = 8'b00010010;
		color_arr[10624] = 8'b00010010;
		color_arr[10625] = 8'b00000000;
		color_arr[10626] = 8'b00000000;
		color_arr[10627] = 8'b00010010;
		color_arr[10628] = 8'b00010010;
		color_arr[10629] = 8'b00010010;
		color_arr[10630] = 8'b00010010;
		color_arr[10631] = 8'b00010010;
		color_arr[10632] = 8'b00010010;
		color_arr[10633] = 8'b00010010;
		color_arr[10634] = 8'b00010010;
		color_arr[10635] = 8'b00010010;
		color_arr[10636] = 8'b00010010;
		color_arr[10637] = 8'b00010010;
		color_arr[10638] = 8'b00010010;
		color_arr[10639] = 8'b00010010;
		color_arr[10640] = 8'b00010010;
		color_arr[10641] = 8'b00010010;
		color_arr[10642] = 8'b00100000;
		color_arr[10643] = 8'b00100000;
		color_arr[10644] = 8'b00100000;
		color_arr[10645] = 8'b00100000;
		color_arr[10646] = 8'b00000000;
		color_arr[10647] = 8'b00000000;
		color_arr[10648] = 8'b00100000;
		color_arr[10649] = 8'b00100000;
		color_arr[10650] = 8'b00100000;
		color_arr[10651] = 8'b00100000;
		color_arr[10652] = 8'b00100000;
		color_arr[10653] = 8'b00100000;
		color_arr[10654] = 8'b00100000;
		color_arr[10655] = 8'b00100000;
		color_arr[10656] = 8'b00100000;
		color_arr[10657] = 8'b00100000;
		color_arr[10658] = 8'b00100000;
		color_arr[10659] = 8'b00100000;
		color_arr[10660] = 8'b00100000;
		color_arr[10661] = 8'b00100000;
		color_arr[10662] = 8'b00100000;
		color_arr[10663] = 8'b00100000;
		color_arr[10664] = 8'b00100000;
		color_arr[10665] = 8'b00100000;
		color_arr[10666] = 8'b00100000;
		color_arr[10667] = 8'b00100000;
		color_arr[10668] = 8'b00100000;
		color_arr[10669] = 8'b00100000;
		color_arr[10670] = 8'b00100000;
		color_arr[10671] = 8'b00100000;
		color_arr[10672] = 8'b00100000;
		color_arr[10673] = 8'b00100000;
		color_arr[10674] = 8'b00100000;
		color_arr[10675] = 8'b00100000;
		color_arr[10676] = 8'b00100000;
		color_arr[10677] = 8'b00100000;
		color_arr[10678] = 8'b00100000;
		color_arr[10679] = 8'b00100000;
		color_arr[10680] = 8'b00100000;
		color_arr[10681] = 8'b00100000;
		color_arr[10682] = 8'b00100000;
		color_arr[10683] = 8'b00100000;
		color_arr[10684] = 8'b00100000;
		color_arr[10685] = 8'b00100000;
		color_arr[10686] = 8'b00100000;
		color_arr[10687] = 8'b00100000;
		color_arr[10688] = 8'b00100000;
		color_arr[10689] = 8'b00100000;
		color_arr[10690] = 8'b00100000;
		color_arr[10691] = 8'b00100000;
		color_arr[10692] = 8'b00100000;
		color_arr[10693] = 8'b00100000;
		color_arr[10694] = 8'b00100000;
		color_arr[10695] = 8'b00100000;
		color_arr[10696] = 8'b00100000;
		color_arr[10697] = 8'b00100000;
		color_arr[10698] = 8'b00100000;
		color_arr[10699] = 8'b00100000;
		color_arr[10700] = 8'b00100000;
		color_arr[10701] = 8'b00000000;
		color_arr[10702] = 8'b00000000;
		color_arr[10703] = 8'b00000000;
		color_arr[10704] = 8'b00001000;
		color_arr[10705] = 8'b00001000;
		color_arr[10706] = 8'b00001000;
		color_arr[10707] = 8'b00001000;
		color_arr[10708] = 8'b00001000;
		color_arr[10709] = 8'b00001000;
		color_arr[10710] = 8'b00001000;
		color_arr[10711] = 8'b00001000;
		color_arr[10712] = 8'b00001000;
		color_arr[10713] = 8'b00001000;
		color_arr[10714] = 8'b00001000;
		color_arr[10715] = 8'b00001000;
		color_arr[10716] = 8'b00001000;
		color_arr[10717] = 8'b00001000;
		color_arr[10718] = 8'b00001000;
		color_arr[10719] = 8'b00001000;
		color_arr[10720] = 8'b00001000;
		color_arr[10721] = 8'b00001000;
		color_arr[10722] = 8'b00001000;
		color_arr[10723] = 8'b00001000;
		color_arr[10724] = 8'b00001000;
		color_arr[10725] = 8'b00001000;
		color_arr[10726] = 8'b00001000;
		color_arr[10727] = 8'b00001000;
		color_arr[10728] = 8'b00001000;
		color_arr[10729] = 8'b00001000;
		color_arr[10730] = 8'b00001000;
		color_arr[10731] = 8'b00001000;
		color_arr[10732] = 8'b00001000;
		color_arr[10733] = 8'b00001000;
		color_arr[10734] = 8'b00001000;
		color_arr[10735] = 8'b00001000;
		color_arr[10736] = 8'b00001000;
		color_arr[10737] = 8'b00001000;
		color_arr[10738] = 8'b00001000;
		color_arr[10739] = 8'b00001000;
		color_arr[10740] = 8'b00001000;
		color_arr[10741] = 8'b00000000;
		color_arr[10742] = 8'b00000000;
		color_arr[10743] = 8'b00000000;
		color_arr[10744] = 8'b00000000;
		color_arr[10745] = 8'b00001000;
		color_arr[10746] = 8'b00001000;
		color_arr[10747] = 8'b00001000;
		color_arr[10748] = 8'b00001000;
		color_arr[10749] = 8'b00010010;
		color_arr[10750] = 8'b00010010;
		color_arr[10751] = 8'b00010010;
		color_arr[10752] = 8'b00010010;
		color_arr[10753] = 8'b00000000;
		color_arr[10754] = 8'b00000000;
		color_arr[10755] = 8'b00010010;
		color_arr[10756] = 8'b00010010;
		color_arr[10757] = 8'b00010010;
		color_arr[10758] = 8'b00010010;
		color_arr[10759] = 8'b00010010;
		color_arr[10760] = 8'b00010010;
		color_arr[10761] = 8'b00010010;
		color_arr[10762] = 8'b00010010;
		color_arr[10763] = 8'b00010010;
		color_arr[10764] = 8'b00010010;
		color_arr[10765] = 8'b00010010;
		color_arr[10766] = 8'b00010010;
		color_arr[10767] = 8'b00010010;
		color_arr[10768] = 8'b00010010;
		color_arr[10769] = 8'b00010010;
		color_arr[10770] = 8'b00100000;
		color_arr[10771] = 8'b00100000;
		color_arr[10772] = 8'b00100000;
		color_arr[10773] = 8'b00100000;
		color_arr[10774] = 8'b00000000;
		color_arr[10775] = 8'b00000000;
		color_arr[10776] = 8'b00100000;
		color_arr[10777] = 8'b00100000;
		color_arr[10778] = 8'b00100000;
		color_arr[10779] = 8'b00100000;
		color_arr[10780] = 8'b00100000;
		color_arr[10781] = 8'b00100000;
		color_arr[10782] = 8'b00100000;
		color_arr[10783] = 8'b00100000;
		color_arr[10784] = 8'b00100000;
		color_arr[10785] = 8'b00100000;
		color_arr[10786] = 8'b00100000;
		color_arr[10787] = 8'b00100000;
		color_arr[10788] = 8'b00100000;
		color_arr[10789] = 8'b00100000;
		color_arr[10790] = 8'b00100000;
		color_arr[10791] = 8'b00100000;
		color_arr[10792] = 8'b00100000;
		color_arr[10793] = 8'b00100000;
		color_arr[10794] = 8'b00100000;
		color_arr[10795] = 8'b00100000;
		color_arr[10796] = 8'b00100000;
		color_arr[10797] = 8'b00100000;
		color_arr[10798] = 8'b00100000;
		color_arr[10799] = 8'b00100000;
		color_arr[10800] = 8'b00100000;
		color_arr[10801] = 8'b00100000;
		color_arr[10802] = 8'b00100000;
		color_arr[10803] = 8'b00100000;
		color_arr[10804] = 8'b00100000;
		color_arr[10805] = 8'b00100000;
		color_arr[10806] = 8'b00100000;
		color_arr[10807] = 8'b00100000;
		color_arr[10808] = 8'b00100000;
		color_arr[10809] = 8'b00100000;
		color_arr[10810] = 8'b00100000;
		color_arr[10811] = 8'b00100000;
		color_arr[10812] = 8'b00100000;
		color_arr[10813] = 8'b00100000;
		color_arr[10814] = 8'b00100000;
		color_arr[10815] = 8'b00100000;
		color_arr[10816] = 8'b00100000;
		color_arr[10817] = 8'b00100000;
		color_arr[10818] = 8'b00100000;
		color_arr[10819] = 8'b00100000;
		color_arr[10820] = 8'b00100000;
		color_arr[10821] = 8'b00100000;
		color_arr[10822] = 8'b00100000;
		color_arr[10823] = 8'b00100000;
		color_arr[10824] = 8'b00100000;
		color_arr[10825] = 8'b00100000;
		color_arr[10826] = 8'b00100000;
		color_arr[10827] = 8'b00100000;
		color_arr[10828] = 8'b00000000;
		color_arr[10829] = 8'b00000000;
		color_arr[10830] = 8'b00000000;
		color_arr[10831] = 8'b00100000;
		color_arr[10832] = 8'b00001000;
		color_arr[10833] = 8'b00001000;
		color_arr[10834] = 8'b00001000;
		color_arr[10835] = 8'b00001000;
		color_arr[10836] = 8'b00001000;
		color_arr[10837] = 8'b00001000;
		color_arr[10838] = 8'b00001000;
		color_arr[10839] = 8'b00001000;
		color_arr[10840] = 8'b00001000;
		color_arr[10841] = 8'b00001000;
		color_arr[10842] = 8'b00001000;
		color_arr[10843] = 8'b00001000;
		color_arr[10844] = 8'b00001000;
		color_arr[10845] = 8'b00001000;
		color_arr[10846] = 8'b00001000;
		color_arr[10847] = 8'b00001000;
		color_arr[10848] = 8'b00001000;
		color_arr[10849] = 8'b00001000;
		color_arr[10850] = 8'b00001000;
		color_arr[10851] = 8'b00001000;
		color_arr[10852] = 8'b00001000;
		color_arr[10853] = 8'b00001000;
		color_arr[10854] = 8'b00001000;
		color_arr[10855] = 8'b00001000;
		color_arr[10856] = 8'b00001000;
		color_arr[10857] = 8'b00001000;
		color_arr[10858] = 8'b00001000;
		color_arr[10859] = 8'b00001000;
		color_arr[10860] = 8'b00001000;
		color_arr[10861] = 8'b00001000;
		color_arr[10862] = 8'b00001000;
		color_arr[10863] = 8'b00001000;
		color_arr[10864] = 8'b00001000;
		color_arr[10865] = 8'b00001000;
		color_arr[10866] = 8'b00001000;
		color_arr[10867] = 8'b00001000;
		color_arr[10868] = 8'b00001000;
		color_arr[10869] = 8'b00000000;
		color_arr[10870] = 8'b00000000;
		color_arr[10871] = 8'b00000000;
		color_arr[10872] = 8'b00000000;
		color_arr[10873] = 8'b00001000;
		color_arr[10874] = 8'b00001000;
		color_arr[10875] = 8'b00001000;
		color_arr[10876] = 8'b00001000;
		color_arr[10877] = 8'b00010010;
		color_arr[10878] = 8'b00010010;
		color_arr[10879] = 8'b00010010;
		color_arr[10880] = 8'b00000000;
		color_arr[10881] = 8'b00000000;
		color_arr[10882] = 8'b00000000;
		color_arr[10883] = 8'b00010010;
		color_arr[10884] = 8'b00010010;
		color_arr[10885] = 8'b00010010;
		color_arr[10886] = 8'b00010010;
		color_arr[10887] = 8'b00010010;
		color_arr[10888] = 8'b00010010;
		color_arr[10889] = 8'b00010010;
		color_arr[10890] = 8'b00010010;
		color_arr[10891] = 8'b00010010;
		color_arr[10892] = 8'b00010010;
		color_arr[10893] = 8'b00010010;
		color_arr[10894] = 8'b00010010;
		color_arr[10895] = 8'b00010010;
		color_arr[10896] = 8'b00010010;
		color_arr[10897] = 8'b00010010;
		color_arr[10898] = 8'b00100000;
		color_arr[10899] = 8'b00100000;
		color_arr[10900] = 8'b00100000;
		color_arr[10901] = 8'b00100000;
		color_arr[10902] = 8'b00000000;
		color_arr[10903] = 8'b00000000;
		color_arr[10904] = 8'b00100000;
		color_arr[10905] = 8'b00100000;
		color_arr[10906] = 8'b00100000;
		color_arr[10907] = 8'b00100000;
		color_arr[10908] = 8'b00100000;
		color_arr[10909] = 8'b00100000;
		color_arr[10910] = 8'b00100000;
		color_arr[10911] = 8'b00100000;
		color_arr[10912] = 8'b00100000;
		color_arr[10913] = 8'b00100000;
		color_arr[10914] = 8'b00100000;
		color_arr[10915] = 8'b00100000;
		color_arr[10916] = 8'b00100000;
		color_arr[10917] = 8'b00100000;
		color_arr[10918] = 8'b00100000;
		color_arr[10919] = 8'b00100000;
		color_arr[10920] = 8'b00100000;
		color_arr[10921] = 8'b00100000;
		color_arr[10922] = 8'b00100000;
		color_arr[10923] = 8'b00100000;
		color_arr[10924] = 8'b00100000;
		color_arr[10925] = 8'b00100000;
		color_arr[10926] = 8'b00100000;
		color_arr[10927] = 8'b00100000;
		color_arr[10928] = 8'b00100000;
		color_arr[10929] = 8'b00100000;
		color_arr[10930] = 8'b00100000;
		color_arr[10931] = 8'b00100000;
		color_arr[10932] = 8'b00100000;
		color_arr[10933] = 8'b00100000;
		color_arr[10934] = 8'b00100000;
		color_arr[10935] = 8'b00100000;
		color_arr[10936] = 8'b00100000;
		color_arr[10937] = 8'b00100000;
		color_arr[10938] = 8'b00100000;
		color_arr[10939] = 8'b00100000;
		color_arr[10940] = 8'b00100000;
		color_arr[10941] = 8'b00100000;
		color_arr[10942] = 8'b00100000;
		color_arr[10943] = 8'b00100000;
		color_arr[10944] = 8'b00100000;
		color_arr[10945] = 8'b00100000;
		color_arr[10946] = 8'b00100000;
		color_arr[10947] = 8'b00100000;
		color_arr[10948] = 8'b00100000;
		color_arr[10949] = 8'b00100000;
		color_arr[10950] = 8'b00100000;
		color_arr[10951] = 8'b00100000;
		color_arr[10952] = 8'b00100000;
		color_arr[10953] = 8'b00100000;
		color_arr[10954] = 8'b00100000;
		color_arr[10955] = 8'b00000000;
		color_arr[10956] = 8'b00000000;
		color_arr[10957] = 8'b00000000;
		color_arr[10958] = 8'b00100000;
		color_arr[10959] = 8'b00100000;
		color_arr[10960] = 8'b00001000;
		color_arr[10961] = 8'b00001000;
		color_arr[10962] = 8'b00001000;
		color_arr[10963] = 8'b00001000;
		color_arr[10964] = 8'b00001000;
		color_arr[10965] = 8'b00001000;
		color_arr[10966] = 8'b00001000;
		color_arr[10967] = 8'b00001000;
		color_arr[10968] = 8'b00001000;
		color_arr[10969] = 8'b00001000;
		color_arr[10970] = 8'b00001000;
		color_arr[10971] = 8'b00001000;
		color_arr[10972] = 8'b00001000;
		color_arr[10973] = 8'b00001000;
		color_arr[10974] = 8'b00001000;
		color_arr[10975] = 8'b00001000;
		color_arr[10976] = 8'b00001000;
		color_arr[10977] = 8'b00001000;
		color_arr[10978] = 8'b00001000;
		color_arr[10979] = 8'b00001000;
		color_arr[10980] = 8'b00001000;
		color_arr[10981] = 8'b00001000;
		color_arr[10982] = 8'b00001000;
		color_arr[10983] = 8'b00001000;
		color_arr[10984] = 8'b00001000;
		color_arr[10985] = 8'b00001000;
		color_arr[10986] = 8'b00001000;
		color_arr[10987] = 8'b00001000;
		color_arr[10988] = 8'b00001000;
		color_arr[10989] = 8'b00001000;
		color_arr[10990] = 8'b00001000;
		color_arr[10991] = 8'b00001000;
		color_arr[10992] = 8'b00001000;
		color_arr[10993] = 8'b00001000;
		color_arr[10994] = 8'b00001000;
		color_arr[10995] = 8'b00001000;
		color_arr[10996] = 8'b00001000;
		color_arr[10997] = 8'b00000000;
		color_arr[10998] = 8'b00000000;
		color_arr[10999] = 8'b00000000;
		color_arr[11000] = 8'b00000000;
		color_arr[11001] = 8'b00001000;
		color_arr[11002] = 8'b00001000;
		color_arr[11003] = 8'b00001000;
		color_arr[11004] = 8'b00001000;
		color_arr[11005] = 8'b00010010;
		color_arr[11006] = 8'b00010010;
		color_arr[11007] = 8'b00010010;
		color_arr[11008] = 8'b00000000;
		color_arr[11009] = 8'b00000000;
		color_arr[11010] = 8'b00010010;
		color_arr[11011] = 8'b00010010;
		color_arr[11012] = 8'b00010010;
		color_arr[11013] = 8'b00010010;
		color_arr[11014] = 8'b00010010;
		color_arr[11015] = 8'b00010010;
		color_arr[11016] = 8'b00010010;
		color_arr[11017] = 8'b00010010;
		color_arr[11018] = 8'b00010010;
		color_arr[11019] = 8'b00010010;
		color_arr[11020] = 8'b00010010;
		color_arr[11021] = 8'b00010010;
		color_arr[11022] = 8'b00010010;
		color_arr[11023] = 8'b00010010;
		color_arr[11024] = 8'b00010010;
		color_arr[11025] = 8'b00010010;
		color_arr[11026] = 8'b00100000;
		color_arr[11027] = 8'b00100000;
		color_arr[11028] = 8'b00100000;
		color_arr[11029] = 8'b00100000;
		color_arr[11030] = 8'b00000000;
		color_arr[11031] = 8'b00000000;
		color_arr[11032] = 8'b00100000;
		color_arr[11033] = 8'b00100000;
		color_arr[11034] = 8'b00100000;
		color_arr[11035] = 8'b00100000;
		color_arr[11036] = 8'b00100000;
		color_arr[11037] = 8'b00100000;
		color_arr[11038] = 8'b00100000;
		color_arr[11039] = 8'b00100000;
		color_arr[11040] = 8'b00100000;
		color_arr[11041] = 8'b00100000;
		color_arr[11042] = 8'b00100000;
		color_arr[11043] = 8'b00100000;
		color_arr[11044] = 8'b00100000;
		color_arr[11045] = 8'b00100000;
		color_arr[11046] = 8'b00100000;
		color_arr[11047] = 8'b00100000;
		color_arr[11048] = 8'b00100000;
		color_arr[11049] = 8'b00100000;
		color_arr[11050] = 8'b00100000;
		color_arr[11051] = 8'b00100000;
		color_arr[11052] = 8'b00100000;
		color_arr[11053] = 8'b00100000;
		color_arr[11054] = 8'b00100000;
		color_arr[11055] = 8'b00100000;
		color_arr[11056] = 8'b00100000;
		color_arr[11057] = 8'b00100000;
		color_arr[11058] = 8'b00100000;
		color_arr[11059] = 8'b00100000;
		color_arr[11060] = 8'b00100000;
		color_arr[11061] = 8'b00100000;
		color_arr[11062] = 8'b00100000;
		color_arr[11063] = 8'b00100000;
		color_arr[11064] = 8'b00100000;
		color_arr[11065] = 8'b00100000;
		color_arr[11066] = 8'b00100000;
		color_arr[11067] = 8'b00100000;
		color_arr[11068] = 8'b00100000;
		color_arr[11069] = 8'b00100000;
		color_arr[11070] = 8'b00100000;
		color_arr[11071] = 8'b00100000;
		color_arr[11072] = 8'b00100000;
		color_arr[11073] = 8'b00100000;
		color_arr[11074] = 8'b00100000;
		color_arr[11075] = 8'b00100000;
		color_arr[11076] = 8'b00100000;
		color_arr[11077] = 8'b00100000;
		color_arr[11078] = 8'b00100000;
		color_arr[11079] = 8'b00100000;
		color_arr[11080] = 8'b00100000;
		color_arr[11081] = 8'b00000000;
		color_arr[11082] = 8'b00000000;
		color_arr[11083] = 8'b00000000;
		color_arr[11084] = 8'b00000000;
		color_arr[11085] = 8'b00100000;
		color_arr[11086] = 8'b00100000;
		color_arr[11087] = 8'b00100000;
		color_arr[11088] = 8'b00001000;
		color_arr[11089] = 8'b00001000;
		color_arr[11090] = 8'b00001000;
		color_arr[11091] = 8'b00001000;
		color_arr[11092] = 8'b00001000;
		color_arr[11093] = 8'b00001000;
		color_arr[11094] = 8'b00001000;
		color_arr[11095] = 8'b00001000;
		color_arr[11096] = 8'b00001000;
		color_arr[11097] = 8'b00001000;
		color_arr[11098] = 8'b00001000;
		color_arr[11099] = 8'b00001000;
		color_arr[11100] = 8'b00001000;
		color_arr[11101] = 8'b00001000;
		color_arr[11102] = 8'b00001000;
		color_arr[11103] = 8'b00001000;
		color_arr[11104] = 8'b00001000;
		color_arr[11105] = 8'b00001000;
		color_arr[11106] = 8'b00001000;
		color_arr[11107] = 8'b00001000;
		color_arr[11108] = 8'b00001000;
		color_arr[11109] = 8'b00001000;
		color_arr[11110] = 8'b00001000;
		color_arr[11111] = 8'b00001000;
		color_arr[11112] = 8'b00001000;
		color_arr[11113] = 8'b00001000;
		color_arr[11114] = 8'b00001000;
		color_arr[11115] = 8'b00001000;
		color_arr[11116] = 8'b00001000;
		color_arr[11117] = 8'b00001000;
		color_arr[11118] = 8'b00001000;
		color_arr[11119] = 8'b00001000;
		color_arr[11120] = 8'b00001000;
		color_arr[11121] = 8'b00001000;
		color_arr[11122] = 8'b00001000;
		color_arr[11123] = 8'b00001000;
		color_arr[11124] = 8'b00000000;
		color_arr[11125] = 8'b00000000;
		color_arr[11126] = 8'b00000000;
		color_arr[11127] = 8'b00000000;
		color_arr[11128] = 8'b00000000;
		color_arr[11129] = 8'b00001000;
		color_arr[11130] = 8'b00001000;
		color_arr[11131] = 8'b00001000;
		color_arr[11132] = 8'b00001000;
		color_arr[11133] = 8'b00010010;
		color_arr[11134] = 8'b00010010;
		color_arr[11135] = 8'b00010010;
		color_arr[11136] = 8'b00000000;
		color_arr[11137] = 8'b00000000;
		color_arr[11138] = 8'b00010010;
		color_arr[11139] = 8'b00010010;
		color_arr[11140] = 8'b00010010;
		color_arr[11141] = 8'b00010010;
		color_arr[11142] = 8'b00010010;
		color_arr[11143] = 8'b00010010;
		color_arr[11144] = 8'b00010010;
		color_arr[11145] = 8'b00010010;
		color_arr[11146] = 8'b00010010;
		color_arr[11147] = 8'b00010010;
		color_arr[11148] = 8'b00010010;
		color_arr[11149] = 8'b00010010;
		color_arr[11150] = 8'b00010010;
		color_arr[11151] = 8'b00010010;
		color_arr[11152] = 8'b00010010;
		color_arr[11153] = 8'b00010010;
		color_arr[11154] = 8'b00100000;
		color_arr[11155] = 8'b00100000;
		color_arr[11156] = 8'b00100000;
		color_arr[11157] = 8'b00100000;
		color_arr[11158] = 8'b00000000;
		color_arr[11159] = 8'b00000000;
		color_arr[11160] = 8'b00100000;
		color_arr[11161] = 8'b00100000;
		color_arr[11162] = 8'b00100000;
		color_arr[11163] = 8'b00100000;
		color_arr[11164] = 8'b00100000;
		color_arr[11165] = 8'b00100000;
		color_arr[11166] = 8'b00100000;
		color_arr[11167] = 8'b00100000;
		color_arr[11168] = 8'b00100000;
		color_arr[11169] = 8'b00100000;
		color_arr[11170] = 8'b00100000;
		color_arr[11171] = 8'b00100000;
		color_arr[11172] = 8'b00100000;
		color_arr[11173] = 8'b00100000;
		color_arr[11174] = 8'b00100000;
		color_arr[11175] = 8'b00100000;
		color_arr[11176] = 8'b00100000;
		color_arr[11177] = 8'b00100000;
		color_arr[11178] = 8'b00100000;
		color_arr[11179] = 8'b00100000;
		color_arr[11180] = 8'b00100000;
		color_arr[11181] = 8'b00100000;
		color_arr[11182] = 8'b00100000;
		color_arr[11183] = 8'b00100000;
		color_arr[11184] = 8'b00100000;
		color_arr[11185] = 8'b00100000;
		color_arr[11186] = 8'b00100000;
		color_arr[11187] = 8'b00100000;
		color_arr[11188] = 8'b00100000;
		color_arr[11189] = 8'b00100000;
		color_arr[11190] = 8'b00100000;
		color_arr[11191] = 8'b00100000;
		color_arr[11192] = 8'b00100000;
		color_arr[11193] = 8'b00100000;
		color_arr[11194] = 8'b00100000;
		color_arr[11195] = 8'b00100000;
		color_arr[11196] = 8'b00100000;
		color_arr[11197] = 8'b00100000;
		color_arr[11198] = 8'b00100000;
		color_arr[11199] = 8'b00100000;
		color_arr[11200] = 8'b00100000;
		color_arr[11201] = 8'b00100000;
		color_arr[11202] = 8'b00100000;
		color_arr[11203] = 8'b00100000;
		color_arr[11204] = 8'b00100000;
		color_arr[11205] = 8'b00100000;
		color_arr[11206] = 8'b00100000;
		color_arr[11207] = 8'b00100000;
		color_arr[11208] = 8'b00000000;
		color_arr[11209] = 8'b00000000;
		color_arr[11210] = 8'b00000000;
		color_arr[11211] = 8'b00000000;
		color_arr[11212] = 8'b00100000;
		color_arr[11213] = 8'b00100000;
		color_arr[11214] = 8'b00100000;
		color_arr[11215] = 8'b00100000;
		color_arr[11216] = 8'b00001000;
		color_arr[11217] = 8'b00001000;
		color_arr[11218] = 8'b00001000;
		color_arr[11219] = 8'b00001000;
		color_arr[11220] = 8'b00001000;
		color_arr[11221] = 8'b00001000;
		color_arr[11222] = 8'b00001000;
		color_arr[11223] = 8'b00001000;
		color_arr[11224] = 8'b00001000;
		color_arr[11225] = 8'b00001000;
		color_arr[11226] = 8'b00001000;
		color_arr[11227] = 8'b00001000;
		color_arr[11228] = 8'b00001000;
		color_arr[11229] = 8'b00001000;
		color_arr[11230] = 8'b00001000;
		color_arr[11231] = 8'b00001000;
		color_arr[11232] = 8'b00001000;
		color_arr[11233] = 8'b00001000;
		color_arr[11234] = 8'b00001000;
		color_arr[11235] = 8'b00001000;
		color_arr[11236] = 8'b00001000;
		color_arr[11237] = 8'b00001000;
		color_arr[11238] = 8'b00001000;
		color_arr[11239] = 8'b00001000;
		color_arr[11240] = 8'b00001000;
		color_arr[11241] = 8'b00001000;
		color_arr[11242] = 8'b00001000;
		color_arr[11243] = 8'b00001000;
		color_arr[11244] = 8'b00001000;
		color_arr[11245] = 8'b00001000;
		color_arr[11246] = 8'b00001000;
		color_arr[11247] = 8'b00001000;
		color_arr[11248] = 8'b00001000;
		color_arr[11249] = 8'b00001000;
		color_arr[11250] = 8'b00001000;
		color_arr[11251] = 8'b00001000;
		color_arr[11252] = 8'b00000000;
		color_arr[11253] = 8'b00000000;
		color_arr[11254] = 8'b00001000;
		color_arr[11255] = 8'b00000000;
		color_arr[11256] = 8'b00000000;
		color_arr[11257] = 8'b00001000;
		color_arr[11258] = 8'b00001000;
		color_arr[11259] = 8'b00001000;
		color_arr[11260] = 8'b00001000;
		color_arr[11261] = 8'b00010010;
		color_arr[11262] = 8'b00010010;
		color_arr[11263] = 8'b00010010;
		color_arr[11264] = 8'b00000000;
		color_arr[11265] = 8'b00010010;
		color_arr[11266] = 8'b00010010;
		color_arr[11267] = 8'b00010010;
		color_arr[11268] = 8'b00010010;
		color_arr[11269] = 8'b00010010;
		color_arr[11270] = 8'b00010010;
		color_arr[11271] = 8'b00010010;
		color_arr[11272] = 8'b00010010;
		color_arr[11273] = 8'b00010010;
		color_arr[11274] = 8'b00010010;
		color_arr[11275] = 8'b00010010;
		color_arr[11276] = 8'b00010010;
		color_arr[11277] = 8'b00010010;
		color_arr[11278] = 8'b00010010;
		color_arr[11279] = 8'b00010010;
		color_arr[11280] = 8'b00010010;
		color_arr[11281] = 8'b00010010;
		color_arr[11282] = 8'b00100000;
		color_arr[11283] = 8'b00100000;
		color_arr[11284] = 8'b00100000;
		color_arr[11285] = 8'b00100000;
		color_arr[11286] = 8'b00000000;
		color_arr[11287] = 8'b00000000;
		color_arr[11288] = 8'b00100000;
		color_arr[11289] = 8'b00100000;
		color_arr[11290] = 8'b00100000;
		color_arr[11291] = 8'b00100000;
		color_arr[11292] = 8'b00100000;
		color_arr[11293] = 8'b00100000;
		color_arr[11294] = 8'b00100000;
		color_arr[11295] = 8'b00100000;
		color_arr[11296] = 8'b00100000;
		color_arr[11297] = 8'b00100000;
		color_arr[11298] = 8'b00100000;
		color_arr[11299] = 8'b00100000;
		color_arr[11300] = 8'b00100000;
		color_arr[11301] = 8'b00100000;
		color_arr[11302] = 8'b00100000;
		color_arr[11303] = 8'b00100000;
		color_arr[11304] = 8'b00100000;
		color_arr[11305] = 8'b00100000;
		color_arr[11306] = 8'b00100000;
		color_arr[11307] = 8'b00100000;
		color_arr[11308] = 8'b00100000;
		color_arr[11309] = 8'b00100000;
		color_arr[11310] = 8'b00100000;
		color_arr[11311] = 8'b00100000;
		color_arr[11312] = 8'b00100000;
		color_arr[11313] = 8'b00100000;
		color_arr[11314] = 8'b00100000;
		color_arr[11315] = 8'b00100000;
		color_arr[11316] = 8'b00100000;
		color_arr[11317] = 8'b00100000;
		color_arr[11318] = 8'b00100000;
		color_arr[11319] = 8'b00100000;
		color_arr[11320] = 8'b00100000;
		color_arr[11321] = 8'b00100000;
		color_arr[11322] = 8'b00100000;
		color_arr[11323] = 8'b00100000;
		color_arr[11324] = 8'b00100000;
		color_arr[11325] = 8'b00100000;
		color_arr[11326] = 8'b00100000;
		color_arr[11327] = 8'b00100000;
		color_arr[11328] = 8'b00100000;
		color_arr[11329] = 8'b00100000;
		color_arr[11330] = 8'b00100000;
		color_arr[11331] = 8'b00100000;
		color_arr[11332] = 8'b00100000;
		color_arr[11333] = 8'b00100000;
		color_arr[11334] = 8'b00100000;
		color_arr[11335] = 8'b00000000;
		color_arr[11336] = 8'b00000000;
		color_arr[11337] = 8'b00000000;
		color_arr[11338] = 8'b00100000;
		color_arr[11339] = 8'b00100000;
		color_arr[11340] = 8'b00100000;
		color_arr[11341] = 8'b00100000;
		color_arr[11342] = 8'b00100000;
		color_arr[11343] = 8'b00100000;
		color_arr[11344] = 8'b00001000;
		color_arr[11345] = 8'b00001000;
		color_arr[11346] = 8'b00001000;
		color_arr[11347] = 8'b00001000;
		color_arr[11348] = 8'b00001000;
		color_arr[11349] = 8'b00001000;
		color_arr[11350] = 8'b00001000;
		color_arr[11351] = 8'b00001000;
		color_arr[11352] = 8'b00001000;
		color_arr[11353] = 8'b00001000;
		color_arr[11354] = 8'b00001000;
		color_arr[11355] = 8'b00001000;
		color_arr[11356] = 8'b00001000;
		color_arr[11357] = 8'b00001000;
		color_arr[11358] = 8'b00001000;
		color_arr[11359] = 8'b00001000;
		color_arr[11360] = 8'b00001000;
		color_arr[11361] = 8'b00001000;
		color_arr[11362] = 8'b00001000;
		color_arr[11363] = 8'b00001000;
		color_arr[11364] = 8'b00001000;
		color_arr[11365] = 8'b00001000;
		color_arr[11366] = 8'b00001000;
		color_arr[11367] = 8'b00001000;
		color_arr[11368] = 8'b00001000;
		color_arr[11369] = 8'b00001000;
		color_arr[11370] = 8'b00001000;
		color_arr[11371] = 8'b00001000;
		color_arr[11372] = 8'b00001000;
		color_arr[11373] = 8'b00001000;
		color_arr[11374] = 8'b00001000;
		color_arr[11375] = 8'b00001000;
		color_arr[11376] = 8'b00001000;
		color_arr[11377] = 8'b00001000;
		color_arr[11378] = 8'b00001000;
		color_arr[11379] = 8'b00001000;
		color_arr[11380] = 8'b00000000;
		color_arr[11381] = 8'b00000000;
		color_arr[11382] = 8'b00001000;
		color_arr[11383] = 8'b00000000;
		color_arr[11384] = 8'b00000000;
		color_arr[11385] = 8'b00001000;
		color_arr[11386] = 8'b00001000;
		color_arr[11387] = 8'b00001000;
		color_arr[11388] = 8'b00001000;
		color_arr[11389] = 8'b00010010;
		color_arr[11390] = 8'b00010010;
		color_arr[11391] = 8'b00010010;
		color_arr[11392] = 8'b00000000;
		color_arr[11393] = 8'b00010010;
		color_arr[11394] = 8'b00010010;
		color_arr[11395] = 8'b00010010;
		color_arr[11396] = 8'b00010010;
		color_arr[11397] = 8'b00010010;
		color_arr[11398] = 8'b00010010;
		color_arr[11399] = 8'b00010010;
		color_arr[11400] = 8'b00010010;
		color_arr[11401] = 8'b00010010;
		color_arr[11402] = 8'b00010010;
		color_arr[11403] = 8'b00010010;
		color_arr[11404] = 8'b00010010;
		color_arr[11405] = 8'b00010010;
		color_arr[11406] = 8'b00010010;
		color_arr[11407] = 8'b00010010;
		color_arr[11408] = 8'b00010010;
		color_arr[11409] = 8'b00010010;
		color_arr[11410] = 8'b00100000;
		color_arr[11411] = 8'b00100000;
		color_arr[11412] = 8'b00100000;
		color_arr[11413] = 8'b00100000;
		color_arr[11414] = 8'b00000000;
		color_arr[11415] = 8'b00000000;
		color_arr[11416] = 8'b00100000;
		color_arr[11417] = 8'b00100000;
		color_arr[11418] = 8'b00100000;
		color_arr[11419] = 8'b00100000;
		color_arr[11420] = 8'b00100000;
		color_arr[11421] = 8'b00100000;
		color_arr[11422] = 8'b00100000;
		color_arr[11423] = 8'b00100000;
		color_arr[11424] = 8'b00100000;
		color_arr[11425] = 8'b00100000;
		color_arr[11426] = 8'b00100000;
		color_arr[11427] = 8'b00100000;
		color_arr[11428] = 8'b00100000;
		color_arr[11429] = 8'b00100000;
		color_arr[11430] = 8'b00100000;
		color_arr[11431] = 8'b00100000;
		color_arr[11432] = 8'b00100000;
		color_arr[11433] = 8'b00100000;
		color_arr[11434] = 8'b00100000;
		color_arr[11435] = 8'b00100000;
		color_arr[11436] = 8'b00100000;
		color_arr[11437] = 8'b00100000;
		color_arr[11438] = 8'b00100000;
		color_arr[11439] = 8'b00100000;
		color_arr[11440] = 8'b00000000;
		color_arr[11441] = 8'b00000000;
		color_arr[11442] = 8'b00000000;
		color_arr[11443] = 8'b00100000;
		color_arr[11444] = 8'b00100000;
		color_arr[11445] = 8'b00100000;
		color_arr[11446] = 8'b00100000;
		color_arr[11447] = 8'b00100000;
		color_arr[11448] = 8'b00100000;
		color_arr[11449] = 8'b00100000;
		color_arr[11450] = 8'b00100000;
		color_arr[11451] = 8'b00100000;
		color_arr[11452] = 8'b00100000;
		color_arr[11453] = 8'b00100000;
		color_arr[11454] = 8'b00100000;
		color_arr[11455] = 8'b00100000;
		color_arr[11456] = 8'b00100000;
		color_arr[11457] = 8'b00100000;
		color_arr[11458] = 8'b00100000;
		color_arr[11459] = 8'b00100000;
		color_arr[11460] = 8'b00100000;
		color_arr[11461] = 8'b00100000;
		color_arr[11462] = 8'b00000000;
		color_arr[11463] = 8'b00000000;
		color_arr[11464] = 8'b00000000;
		color_arr[11465] = 8'b00100000;
		color_arr[11466] = 8'b00100000;
		color_arr[11467] = 8'b00100000;
		color_arr[11468] = 8'b00100000;
		color_arr[11469] = 8'b00100000;
		color_arr[11470] = 8'b00100000;
		color_arr[11471] = 8'b00100000;
		color_arr[11472] = 8'b00001000;
		color_arr[11473] = 8'b00001000;
		color_arr[11474] = 8'b00001000;
		color_arr[11475] = 8'b00001000;
		color_arr[11476] = 8'b00001000;
		color_arr[11477] = 8'b00001000;
		color_arr[11478] = 8'b00001000;
		color_arr[11479] = 8'b00001000;
		color_arr[11480] = 8'b00001000;
		color_arr[11481] = 8'b00001000;
		color_arr[11482] = 8'b00001000;
		color_arr[11483] = 8'b00001000;
		color_arr[11484] = 8'b00001000;
		color_arr[11485] = 8'b00001000;
		color_arr[11486] = 8'b00001000;
		color_arr[11487] = 8'b00001000;
		color_arr[11488] = 8'b00001000;
		color_arr[11489] = 8'b00001000;
		color_arr[11490] = 8'b00001000;
		color_arr[11491] = 8'b00001000;
		color_arr[11492] = 8'b00001000;
		color_arr[11493] = 8'b00001000;
		color_arr[11494] = 8'b00001000;
		color_arr[11495] = 8'b00001000;
		color_arr[11496] = 8'b00001000;
		color_arr[11497] = 8'b00001000;
		color_arr[11498] = 8'b00001000;
		color_arr[11499] = 8'b00001000;
		color_arr[11500] = 8'b00001000;
		color_arr[11501] = 8'b00001000;
		color_arr[11502] = 8'b00001000;
		color_arr[11503] = 8'b00001000;
		color_arr[11504] = 8'b00001000;
		color_arr[11505] = 8'b00001000;
		color_arr[11506] = 8'b00001000;
		color_arr[11507] = 8'b00001000;
		color_arr[11508] = 8'b00000000;
		color_arr[11509] = 8'b00000000;
		color_arr[11510] = 8'b00001000;
		color_arr[11511] = 8'b00000000;
		color_arr[11512] = 8'b00000000;
		color_arr[11513] = 8'b00001000;
		color_arr[11514] = 8'b00001000;
		color_arr[11515] = 8'b00001000;
		color_arr[11516] = 8'b00001000;
		color_arr[11517] = 8'b00010010;
		color_arr[11518] = 8'b00010010;
		color_arr[11519] = 8'b00010010;
		color_arr[11520] = 8'b00000000;
		color_arr[11521] = 8'b00010010;
		color_arr[11522] = 8'b00010010;
		color_arr[11523] = 8'b00010010;
		color_arr[11524] = 8'b00010010;
		color_arr[11525] = 8'b00010010;
		color_arr[11526] = 8'b00010010;
		color_arr[11527] = 8'b00010010;
		color_arr[11528] = 8'b00010010;
		color_arr[11529] = 8'b00010010;
		color_arr[11530] = 8'b00010010;
		color_arr[11531] = 8'b00010010;
		color_arr[11532] = 8'b00010010;
		color_arr[11533] = 8'b00010010;
		color_arr[11534] = 8'b00010010;
		color_arr[11535] = 8'b00010010;
		color_arr[11536] = 8'b00010010;
		color_arr[11537] = 8'b00010010;
		color_arr[11538] = 8'b00100000;
		color_arr[11539] = 8'b00100000;
		color_arr[11540] = 8'b00100000;
		color_arr[11541] = 8'b00100000;
		color_arr[11542] = 8'b00000000;
		color_arr[11543] = 8'b00000000;
		color_arr[11544] = 8'b00100000;
		color_arr[11545] = 8'b00100000;
		color_arr[11546] = 8'b00100000;
		color_arr[11547] = 8'b00100000;
		color_arr[11548] = 8'b00100000;
		color_arr[11549] = 8'b00100000;
		color_arr[11550] = 8'b00100000;
		color_arr[11551] = 8'b00100000;
		color_arr[11552] = 8'b00100000;
		color_arr[11553] = 8'b00100000;
		color_arr[11554] = 8'b00100000;
		color_arr[11555] = 8'b00100000;
		color_arr[11556] = 8'b00100000;
		color_arr[11557] = 8'b00100000;
		color_arr[11558] = 8'b00100000;
		color_arr[11559] = 8'b00100000;
		color_arr[11560] = 8'b00100000;
		color_arr[11561] = 8'b00100000;
		color_arr[11562] = 8'b00100000;
		color_arr[11563] = 8'b00100000;
		color_arr[11564] = 8'b00100000;
		color_arr[11565] = 8'b00100000;
		color_arr[11566] = 8'b00100000;
		color_arr[11567] = 8'b00000000;
		color_arr[11568] = 8'b00000000;
		color_arr[11569] = 8'b00000000;
		color_arr[11570] = 8'b00000000;
		color_arr[11571] = 8'b00100000;
		color_arr[11572] = 8'b00100000;
		color_arr[11573] = 8'b00100000;
		color_arr[11574] = 8'b00100000;
		color_arr[11575] = 8'b00100000;
		color_arr[11576] = 8'b00100000;
		color_arr[11577] = 8'b00100000;
		color_arr[11578] = 8'b00100000;
		color_arr[11579] = 8'b00100000;
		color_arr[11580] = 8'b00100000;
		color_arr[11581] = 8'b00100000;
		color_arr[11582] = 8'b00100000;
		color_arr[11583] = 8'b00100000;
		color_arr[11584] = 8'b00100000;
		color_arr[11585] = 8'b00100000;
		color_arr[11586] = 8'b00100000;
		color_arr[11587] = 8'b00100000;
		color_arr[11588] = 8'b00100000;
		color_arr[11589] = 8'b00000000;
		color_arr[11590] = 8'b00000000;
		color_arr[11591] = 8'b00000000;
		color_arr[11592] = 8'b00100000;
		color_arr[11593] = 8'b00100000;
		color_arr[11594] = 8'b00100000;
		color_arr[11595] = 8'b00100000;
		color_arr[11596] = 8'b00100000;
		color_arr[11597] = 8'b00100000;
		color_arr[11598] = 8'b00100000;
		color_arr[11599] = 8'b00100000;
		color_arr[11600] = 8'b00001000;
		color_arr[11601] = 8'b00001000;
		color_arr[11602] = 8'b00001000;
		color_arr[11603] = 8'b00001000;
		color_arr[11604] = 8'b00001000;
		color_arr[11605] = 8'b00001000;
		color_arr[11606] = 8'b00001000;
		color_arr[11607] = 8'b00001000;
		color_arr[11608] = 8'b00001000;
		color_arr[11609] = 8'b00001000;
		color_arr[11610] = 8'b00001000;
		color_arr[11611] = 8'b00001000;
		color_arr[11612] = 8'b00001000;
		color_arr[11613] = 8'b00001000;
		color_arr[11614] = 8'b00001000;
		color_arr[11615] = 8'b00001000;
		color_arr[11616] = 8'b00001000;
		color_arr[11617] = 8'b00001000;
		color_arr[11618] = 8'b00001000;
		color_arr[11619] = 8'b00001000;
		color_arr[11620] = 8'b00001000;
		color_arr[11621] = 8'b00001000;
		color_arr[11622] = 8'b00001000;
		color_arr[11623] = 8'b00001000;
		color_arr[11624] = 8'b00001000;
		color_arr[11625] = 8'b00001000;
		color_arr[11626] = 8'b00001000;
		color_arr[11627] = 8'b00001000;
		color_arr[11628] = 8'b00001000;
		color_arr[11629] = 8'b00001000;
		color_arr[11630] = 8'b00001000;
		color_arr[11631] = 8'b00001000;
		color_arr[11632] = 8'b00001000;
		color_arr[11633] = 8'b00001000;
		color_arr[11634] = 8'b00001000;
		color_arr[11635] = 8'b00000000;
		color_arr[11636] = 8'b00000000;
		color_arr[11637] = 8'b00000000;
		color_arr[11638] = 8'b00001000;
		color_arr[11639] = 8'b00000000;
		color_arr[11640] = 8'b00000000;
		color_arr[11641] = 8'b00001000;
		color_arr[11642] = 8'b00001000;
		color_arr[11643] = 8'b00001000;
		color_arr[11644] = 8'b00001000;
		color_arr[11645] = 8'b00010010;
		color_arr[11646] = 8'b00010010;
		color_arr[11647] = 8'b00010010;
		color_arr[11648] = 8'b00010010;
		color_arr[11649] = 8'b00010010;
		color_arr[11650] = 8'b00010010;
		color_arr[11651] = 8'b00010010;
		color_arr[11652] = 8'b00010010;
		color_arr[11653] = 8'b00010010;
		color_arr[11654] = 8'b00010010;
		color_arr[11655] = 8'b00010010;
		color_arr[11656] = 8'b00010010;
		color_arr[11657] = 8'b00010010;
		color_arr[11658] = 8'b00010010;
		color_arr[11659] = 8'b00010010;
		color_arr[11660] = 8'b00010010;
		color_arr[11661] = 8'b00010010;
		color_arr[11662] = 8'b00010010;
		color_arr[11663] = 8'b00010010;
		color_arr[11664] = 8'b00010010;
		color_arr[11665] = 8'b00010010;
		color_arr[11666] = 8'b00100000;
		color_arr[11667] = 8'b00100000;
		color_arr[11668] = 8'b00100000;
		color_arr[11669] = 8'b00100000;
		color_arr[11670] = 8'b00000000;
		color_arr[11671] = 8'b00000000;
		color_arr[11672] = 8'b00100000;
		color_arr[11673] = 8'b00100000;
		color_arr[11674] = 8'b00100000;
		color_arr[11675] = 8'b00100000;
		color_arr[11676] = 8'b00100000;
		color_arr[11677] = 8'b00100000;
		color_arr[11678] = 8'b00100000;
		color_arr[11679] = 8'b00100000;
		color_arr[11680] = 8'b00100000;
		color_arr[11681] = 8'b00100000;
		color_arr[11682] = 8'b00100000;
		color_arr[11683] = 8'b00100000;
		color_arr[11684] = 8'b00100000;
		color_arr[11685] = 8'b00100000;
		color_arr[11686] = 8'b00100000;
		color_arr[11687] = 8'b00100000;
		color_arr[11688] = 8'b00100000;
		color_arr[11689] = 8'b00100000;
		color_arr[11690] = 8'b00100000;
		color_arr[11691] = 8'b00100000;
		color_arr[11692] = 8'b00100000;
		color_arr[11693] = 8'b00000000;
		color_arr[11694] = 8'b00000000;
		color_arr[11695] = 8'b00000000;
		color_arr[11696] = 8'b00000000;
		color_arr[11697] = 8'b00100000;
		color_arr[11698] = 8'b00100000;
		color_arr[11699] = 8'b00100000;
		color_arr[11700] = 8'b00100000;
		color_arr[11701] = 8'b00100000;
		color_arr[11702] = 8'b00100000;
		color_arr[11703] = 8'b00100000;
		color_arr[11704] = 8'b00100000;
		color_arr[11705] = 8'b00100000;
		color_arr[11706] = 8'b00100000;
		color_arr[11707] = 8'b00100000;
		color_arr[11708] = 8'b00100000;
		color_arr[11709] = 8'b00100000;
		color_arr[11710] = 8'b00100000;
		color_arr[11711] = 8'b00100000;
		color_arr[11712] = 8'b00100000;
		color_arr[11713] = 8'b00100000;
		color_arr[11714] = 8'b00100000;
		color_arr[11715] = 8'b00000000;
		color_arr[11716] = 8'b00000000;
		color_arr[11717] = 8'b00000000;
		color_arr[11718] = 8'b00000000;
		color_arr[11719] = 8'b00100000;
		color_arr[11720] = 8'b00100000;
		color_arr[11721] = 8'b00100000;
		color_arr[11722] = 8'b00100000;
		color_arr[11723] = 8'b00100000;
		color_arr[11724] = 8'b00100000;
		color_arr[11725] = 8'b00100000;
		color_arr[11726] = 8'b00100000;
		color_arr[11727] = 8'b00100000;
		color_arr[11728] = 8'b00001000;
		color_arr[11729] = 8'b00001000;
		color_arr[11730] = 8'b00001000;
		color_arr[11731] = 8'b00001000;
		color_arr[11732] = 8'b00001000;
		color_arr[11733] = 8'b00001000;
		color_arr[11734] = 8'b00001000;
		color_arr[11735] = 8'b00001000;
		color_arr[11736] = 8'b00001000;
		color_arr[11737] = 8'b00001000;
		color_arr[11738] = 8'b00001000;
		color_arr[11739] = 8'b00001000;
		color_arr[11740] = 8'b00001000;
		color_arr[11741] = 8'b00001000;
		color_arr[11742] = 8'b00001000;
		color_arr[11743] = 8'b00001000;
		color_arr[11744] = 8'b00001000;
		color_arr[11745] = 8'b00001000;
		color_arr[11746] = 8'b00001000;
		color_arr[11747] = 8'b00001000;
		color_arr[11748] = 8'b00001000;
		color_arr[11749] = 8'b00001000;
		color_arr[11750] = 8'b00001000;
		color_arr[11751] = 8'b00001000;
		color_arr[11752] = 8'b00001000;
		color_arr[11753] = 8'b00001000;
		color_arr[11754] = 8'b00001000;
		color_arr[11755] = 8'b00001000;
		color_arr[11756] = 8'b00001000;
		color_arr[11757] = 8'b00001000;
		color_arr[11758] = 8'b00001000;
		color_arr[11759] = 8'b00001000;
		color_arr[11760] = 8'b00001000;
		color_arr[11761] = 8'b00001000;
		color_arr[11762] = 8'b00001000;
		color_arr[11763] = 8'b00000000;
		color_arr[11764] = 8'b00000000;
		color_arr[11765] = 8'b00001000;
		color_arr[11766] = 8'b00001000;
		color_arr[11767] = 8'b00000000;
		color_arr[11768] = 8'b00000000;
		color_arr[11769] = 8'b00001000;
		color_arr[11770] = 8'b00001000;
		color_arr[11771] = 8'b00001000;
		color_arr[11772] = 8'b00001000;
		color_arr[11773] = 8'b00010010;
		color_arr[11774] = 8'b00010010;
		color_arr[11775] = 8'b00010010;
		color_arr[11776] = 8'b00010010;
		color_arr[11777] = 8'b00010010;
		color_arr[11778] = 8'b00010010;
		color_arr[11779] = 8'b00010010;
		color_arr[11780] = 8'b00010010;
		color_arr[11781] = 8'b00010010;
		color_arr[11782] = 8'b00010010;
		color_arr[11783] = 8'b00010010;
		color_arr[11784] = 8'b00010010;
		color_arr[11785] = 8'b00010010;
		color_arr[11786] = 8'b00010010;
		color_arr[11787] = 8'b00010010;
		color_arr[11788] = 8'b00010010;
		color_arr[11789] = 8'b00010010;
		color_arr[11790] = 8'b00010010;
		color_arr[11791] = 8'b00010010;
		color_arr[11792] = 8'b00010010;
		color_arr[11793] = 8'b00010010;
		color_arr[11794] = 8'b00100000;
		color_arr[11795] = 8'b00100000;
		color_arr[11796] = 8'b00100000;
		color_arr[11797] = 8'b00100000;
		color_arr[11798] = 8'b00000000;
		color_arr[11799] = 8'b00000000;
		color_arr[11800] = 8'b00100000;
		color_arr[11801] = 8'b00100000;
		color_arr[11802] = 8'b00100000;
		color_arr[11803] = 8'b00100000;
		color_arr[11804] = 8'b00100000;
		color_arr[11805] = 8'b00100000;
		color_arr[11806] = 8'b00100000;
		color_arr[11807] = 8'b00100000;
		color_arr[11808] = 8'b00100000;
		color_arr[11809] = 8'b00100000;
		color_arr[11810] = 8'b00100000;
		color_arr[11811] = 8'b00100000;
		color_arr[11812] = 8'b00100000;
		color_arr[11813] = 8'b00100000;
		color_arr[11814] = 8'b00100000;
		color_arr[11815] = 8'b00100000;
		color_arr[11816] = 8'b00100000;
		color_arr[11817] = 8'b00100000;
		color_arr[11818] = 8'b00100000;
		color_arr[11819] = 8'b00100000;
		color_arr[11820] = 8'b00000000;
		color_arr[11821] = 8'b00000000;
		color_arr[11822] = 8'b00000000;
		color_arr[11823] = 8'b00000000;
		color_arr[11824] = 8'b00100000;
		color_arr[11825] = 8'b00100000;
		color_arr[11826] = 8'b00100000;
		color_arr[11827] = 8'b00100000;
		color_arr[11828] = 8'b00100000;
		color_arr[11829] = 8'b00100000;
		color_arr[11830] = 8'b00100000;
		color_arr[11831] = 8'b00100000;
		color_arr[11832] = 8'b00100000;
		color_arr[11833] = 8'b00100000;
		color_arr[11834] = 8'b00100000;
		color_arr[11835] = 8'b00100000;
		color_arr[11836] = 8'b00100000;
		color_arr[11837] = 8'b00100000;
		color_arr[11838] = 8'b00100000;
		color_arr[11839] = 8'b00100000;
		color_arr[11840] = 8'b00100000;
		color_arr[11841] = 8'b00100000;
		color_arr[11842] = 8'b00000000;
		color_arr[11843] = 8'b00000000;
		color_arr[11844] = 8'b00000000;
		color_arr[11845] = 8'b00000000;
		color_arr[11846] = 8'b00100000;
		color_arr[11847] = 8'b00100000;
		color_arr[11848] = 8'b00100000;
		color_arr[11849] = 8'b00100000;
		color_arr[11850] = 8'b00100000;
		color_arr[11851] = 8'b00100000;
		color_arr[11852] = 8'b00100000;
		color_arr[11853] = 8'b00100000;
		color_arr[11854] = 8'b00100000;
		color_arr[11855] = 8'b00100000;
		color_arr[11856] = 8'b00001000;
		color_arr[11857] = 8'b00001000;
		color_arr[11858] = 8'b00001000;
		color_arr[11859] = 8'b00001000;
		color_arr[11860] = 8'b00001000;
		color_arr[11861] = 8'b00001000;
		color_arr[11862] = 8'b00001000;
		color_arr[11863] = 8'b00001000;
		color_arr[11864] = 8'b00001000;
		color_arr[11865] = 8'b00001000;
		color_arr[11866] = 8'b00001000;
		color_arr[11867] = 8'b00001000;
		color_arr[11868] = 8'b00001000;
		color_arr[11869] = 8'b00001000;
		color_arr[11870] = 8'b00001000;
		color_arr[11871] = 8'b00001000;
		color_arr[11872] = 8'b00001000;
		color_arr[11873] = 8'b00001000;
		color_arr[11874] = 8'b00001000;
		color_arr[11875] = 8'b00001000;
		color_arr[11876] = 8'b00001000;
		color_arr[11877] = 8'b00001000;
		color_arr[11878] = 8'b00001000;
		color_arr[11879] = 8'b00001000;
		color_arr[11880] = 8'b00001000;
		color_arr[11881] = 8'b00001000;
		color_arr[11882] = 8'b00001000;
		color_arr[11883] = 8'b00001000;
		color_arr[11884] = 8'b00001000;
		color_arr[11885] = 8'b00001000;
		color_arr[11886] = 8'b00001000;
		color_arr[11887] = 8'b00001000;
		color_arr[11888] = 8'b00001000;
		color_arr[11889] = 8'b00001000;
		color_arr[11890] = 8'b00000000;
		color_arr[11891] = 8'b00000000;
		color_arr[11892] = 8'b00000000;
		color_arr[11893] = 8'b00001000;
		color_arr[11894] = 8'b00001000;
		color_arr[11895] = 8'b00000000;
		color_arr[11896] = 8'b00000000;
		color_arr[11897] = 8'b00001000;
		color_arr[11898] = 8'b00001000;
		color_arr[11899] = 8'b00001000;
		color_arr[11900] = 8'b00001000;
		color_arr[11901] = 8'b00010010;
		color_arr[11902] = 8'b00010010;
		color_arr[11903] = 8'b00010010;
		color_arr[11904] = 8'b00010010;
		color_arr[11905] = 8'b00010010;
		color_arr[11906] = 8'b00010010;
		color_arr[11907] = 8'b00010010;
		color_arr[11908] = 8'b00010010;
		color_arr[11909] = 8'b00010010;
		color_arr[11910] = 8'b00010010;
		color_arr[11911] = 8'b00010010;
		color_arr[11912] = 8'b00010010;
		color_arr[11913] = 8'b00010010;
		color_arr[11914] = 8'b00010010;
		color_arr[11915] = 8'b00010010;
		color_arr[11916] = 8'b00010010;
		color_arr[11917] = 8'b00010010;
		color_arr[11918] = 8'b00010010;
		color_arr[11919] = 8'b00010010;
		color_arr[11920] = 8'b00010010;
		color_arr[11921] = 8'b00010010;
		color_arr[11922] = 8'b00100000;
		color_arr[11923] = 8'b00100000;
		color_arr[11924] = 8'b00100000;
		color_arr[11925] = 8'b00100000;
		color_arr[11926] = 8'b00000000;
		color_arr[11927] = 8'b00000000;
		color_arr[11928] = 8'b00100000;
		color_arr[11929] = 8'b00100000;
		color_arr[11930] = 8'b00100000;
		color_arr[11931] = 8'b00100000;
		color_arr[11932] = 8'b00100000;
		color_arr[11933] = 8'b00100000;
		color_arr[11934] = 8'b00100000;
		color_arr[11935] = 8'b00100000;
		color_arr[11936] = 8'b00100000;
		color_arr[11937] = 8'b00100000;
		color_arr[11938] = 8'b00100000;
		color_arr[11939] = 8'b00100000;
		color_arr[11940] = 8'b00100000;
		color_arr[11941] = 8'b00100000;
		color_arr[11942] = 8'b00100000;
		color_arr[11943] = 8'b00100000;
		color_arr[11944] = 8'b00100000;
		color_arr[11945] = 8'b00100000;
		color_arr[11946] = 8'b00000000;
		color_arr[11947] = 8'b00000000;
		color_arr[11948] = 8'b00000000;
		color_arr[11949] = 8'b00000000;
		color_arr[11950] = 8'b00100000;
		color_arr[11951] = 8'b00100000;
		color_arr[11952] = 8'b00100000;
		color_arr[11953] = 8'b00100000;
		color_arr[11954] = 8'b00100000;
		color_arr[11955] = 8'b00100000;
		color_arr[11956] = 8'b00100000;
		color_arr[11957] = 8'b00100000;
		color_arr[11958] = 8'b00100000;
		color_arr[11959] = 8'b00100000;
		color_arr[11960] = 8'b00100000;
		color_arr[11961] = 8'b00100000;
		color_arr[11962] = 8'b00100000;
		color_arr[11963] = 8'b00100000;
		color_arr[11964] = 8'b00100000;
		color_arr[11965] = 8'b00100000;
		color_arr[11966] = 8'b00100000;
		color_arr[11967] = 8'b00100000;
		color_arr[11968] = 8'b00100000;
		color_arr[11969] = 8'b00000000;
		color_arr[11970] = 8'b00000000;
		color_arr[11971] = 8'b00000000;
		color_arr[11972] = 8'b00100000;
		color_arr[11973] = 8'b00100000;
		color_arr[11974] = 8'b00100000;
		color_arr[11975] = 8'b00100000;
		color_arr[11976] = 8'b00100000;
		color_arr[11977] = 8'b00100000;
		color_arr[11978] = 8'b00100000;
		color_arr[11979] = 8'b00100000;
		color_arr[11980] = 8'b00100000;
		color_arr[11981] = 8'b00100000;
		color_arr[11982] = 8'b00100000;
		color_arr[11983] = 8'b00100000;
		color_arr[11984] = 8'b00001000;
		color_arr[11985] = 8'b00001000;
		color_arr[11986] = 8'b00001000;
		color_arr[11987] = 8'b00001000;
		color_arr[11988] = 8'b00001000;
		color_arr[11989] = 8'b00001000;
		color_arr[11990] = 8'b00001000;
		color_arr[11991] = 8'b00001000;
		color_arr[11992] = 8'b00001000;
		color_arr[11993] = 8'b00001000;
		color_arr[11994] = 8'b00001000;
		color_arr[11995] = 8'b00001000;
		color_arr[11996] = 8'b00001000;
		color_arr[11997] = 8'b00001000;
		color_arr[11998] = 8'b00001000;
		color_arr[11999] = 8'b00001000;
		color_arr[12000] = 8'b00001000;
		color_arr[12001] = 8'b00001000;
		color_arr[12002] = 8'b00001000;
		color_arr[12003] = 8'b00001000;
		color_arr[12004] = 8'b00001000;
		color_arr[12005] = 8'b00001000;
		color_arr[12006] = 8'b00001000;
		color_arr[12007] = 8'b00001000;
		color_arr[12008] = 8'b00001000;
		color_arr[12009] = 8'b00001000;
		color_arr[12010] = 8'b00001000;
		color_arr[12011] = 8'b00001000;
		color_arr[12012] = 8'b00001000;
		color_arr[12013] = 8'b00001000;
		color_arr[12014] = 8'b00001000;
		color_arr[12015] = 8'b00001000;
		color_arr[12016] = 8'b00001000;
		color_arr[12017] = 8'b00001000;
		color_arr[12018] = 8'b00000000;
		color_arr[12019] = 8'b00000000;
		color_arr[12020] = 8'b00001000;
		color_arr[12021] = 8'b00001000;
		color_arr[12022] = 8'b00001000;
		color_arr[12023] = 8'b00000000;
		color_arr[12024] = 8'b00000000;
		color_arr[12025] = 8'b00001000;
		color_arr[12026] = 8'b00001000;
		color_arr[12027] = 8'b00001000;
		color_arr[12028] = 8'b00001000;
		color_arr[12029] = 8'b00010010;
		color_arr[12030] = 8'b00010010;
		color_arr[12031] = 8'b00010010;
		color_arr[12032] = 8'b00010010;
		color_arr[12033] = 8'b00010010;
		color_arr[12034] = 8'b00010010;
		color_arr[12035] = 8'b00010010;
		color_arr[12036] = 8'b00010010;
		color_arr[12037] = 8'b00010010;
		color_arr[12038] = 8'b00010010;
		color_arr[12039] = 8'b00010010;
		color_arr[12040] = 8'b00010010;
		color_arr[12041] = 8'b00010010;
		color_arr[12042] = 8'b00010010;
		color_arr[12043] = 8'b00010010;
		color_arr[12044] = 8'b00010010;
		color_arr[12045] = 8'b00010010;
		color_arr[12046] = 8'b00010010;
		color_arr[12047] = 8'b00010010;
		color_arr[12048] = 8'b00010010;
		color_arr[12049] = 8'b00010010;
		color_arr[12050] = 8'b00100000;
		color_arr[12051] = 8'b00100000;
		color_arr[12052] = 8'b00100000;
		color_arr[12053] = 8'b00100000;
		color_arr[12054] = 8'b00000000;
		color_arr[12055] = 8'b00000000;
		color_arr[12056] = 8'b00100000;
		color_arr[12057] = 8'b00100000;
		color_arr[12058] = 8'b00100000;
		color_arr[12059] = 8'b00100000;
		color_arr[12060] = 8'b00100000;
		color_arr[12061] = 8'b00100000;
		color_arr[12062] = 8'b00100000;
		color_arr[12063] = 8'b00100000;
		color_arr[12064] = 8'b00100000;
		color_arr[12065] = 8'b00100000;
		color_arr[12066] = 8'b00100000;
		color_arr[12067] = 8'b00100000;
		color_arr[12068] = 8'b00100000;
		color_arr[12069] = 8'b00100000;
		color_arr[12070] = 8'b00100000;
		color_arr[12071] = 8'b00100000;
		color_arr[12072] = 8'b00100000;
		color_arr[12073] = 8'b00000000;
		color_arr[12074] = 8'b00000000;
		color_arr[12075] = 8'b00000000;
		color_arr[12076] = 8'b00000000;
		color_arr[12077] = 8'b00100000;
		color_arr[12078] = 8'b00100000;
		color_arr[12079] = 8'b00100000;
		color_arr[12080] = 8'b00100000;
		color_arr[12081] = 8'b00100000;
		color_arr[12082] = 8'b00100000;
		color_arr[12083] = 8'b00100000;
		color_arr[12084] = 8'b00100000;
		color_arr[12085] = 8'b00100000;
		color_arr[12086] = 8'b00100000;
		color_arr[12087] = 8'b00100000;
		color_arr[12088] = 8'b00100000;
		color_arr[12089] = 8'b00100000;
		color_arr[12090] = 8'b00100000;
		color_arr[12091] = 8'b00100000;
		color_arr[12092] = 8'b00100000;
		color_arr[12093] = 8'b00100000;
		color_arr[12094] = 8'b00100000;
		color_arr[12095] = 8'b00100000;
		color_arr[12096] = 8'b00000000;
		color_arr[12097] = 8'b00000000;
		color_arr[12098] = 8'b00000000;
		color_arr[12099] = 8'b00100000;
		color_arr[12100] = 8'b00100000;
		color_arr[12101] = 8'b00100000;
		color_arr[12102] = 8'b00100000;
		color_arr[12103] = 8'b00100000;
		color_arr[12104] = 8'b00100000;
		color_arr[12105] = 8'b00100000;
		color_arr[12106] = 8'b00100000;
		color_arr[12107] = 8'b00100000;
		color_arr[12108] = 8'b00100000;
		color_arr[12109] = 8'b00100000;
		color_arr[12110] = 8'b00100000;
		color_arr[12111] = 8'b00100000;
		color_arr[12112] = 8'b00001000;
		color_arr[12113] = 8'b00001000;
		color_arr[12114] = 8'b00001000;
		color_arr[12115] = 8'b00001000;
		color_arr[12116] = 8'b00001000;
		color_arr[12117] = 8'b00001000;
		color_arr[12118] = 8'b00001000;
		color_arr[12119] = 8'b00001000;
		color_arr[12120] = 8'b00001000;
		color_arr[12121] = 8'b00001000;
		color_arr[12122] = 8'b00001000;
		color_arr[12123] = 8'b00001000;
		color_arr[12124] = 8'b00001000;
		color_arr[12125] = 8'b00001000;
		color_arr[12126] = 8'b00001000;
		color_arr[12127] = 8'b00001000;
		color_arr[12128] = 8'b00001000;
		color_arr[12129] = 8'b00001000;
		color_arr[12130] = 8'b00001000;
		color_arr[12131] = 8'b00001000;
		color_arr[12132] = 8'b00001000;
		color_arr[12133] = 8'b00001000;
		color_arr[12134] = 8'b00001000;
		color_arr[12135] = 8'b00001000;
		color_arr[12136] = 8'b00001000;
		color_arr[12137] = 8'b00001000;
		color_arr[12138] = 8'b00001000;
		color_arr[12139] = 8'b00001000;
		color_arr[12140] = 8'b00001000;
		color_arr[12141] = 8'b00001000;
		color_arr[12142] = 8'b00001000;
		color_arr[12143] = 8'b00001000;
		color_arr[12144] = 8'b00001000;
		color_arr[12145] = 8'b00000000;
		color_arr[12146] = 8'b00000000;
		color_arr[12147] = 8'b00000000;
		color_arr[12148] = 8'b00001000;
		color_arr[12149] = 8'b00001000;
		color_arr[12150] = 8'b00001000;
		color_arr[12151] = 8'b00000000;
		color_arr[12152] = 8'b00000000;
		color_arr[12153] = 8'b00001000;
		color_arr[12154] = 8'b00001000;
		color_arr[12155] = 8'b00001000;
		color_arr[12156] = 8'b00001000;
		color_arr[12157] = 8'b00010010;
		color_arr[12158] = 8'b00010010;
		color_arr[12159] = 8'b00010010;
		color_arr[12160] = 8'b00010010;
		color_arr[12161] = 8'b00010010;
		color_arr[12162] = 8'b00010010;
		color_arr[12163] = 8'b00010010;
		color_arr[12164] = 8'b00010010;
		color_arr[12165] = 8'b00010010;
		color_arr[12166] = 8'b00010010;
		color_arr[12167] = 8'b00010010;
		color_arr[12168] = 8'b00010010;
		color_arr[12169] = 8'b00010010;
		color_arr[12170] = 8'b00010010;
		color_arr[12171] = 8'b00010010;
		color_arr[12172] = 8'b00010010;
		color_arr[12173] = 8'b00010010;
		color_arr[12174] = 8'b00010010;
		color_arr[12175] = 8'b00010010;
		color_arr[12176] = 8'b00010010;
		color_arr[12177] = 8'b00010010;
		color_arr[12178] = 8'b00100000;
		color_arr[12179] = 8'b00100000;
		color_arr[12180] = 8'b00100000;
		color_arr[12181] = 8'b00100000;
		color_arr[12182] = 8'b00000000;
		color_arr[12183] = 8'b00000000;
		color_arr[12184] = 8'b00100000;
		color_arr[12185] = 8'b00100000;
		color_arr[12186] = 8'b00100000;
		color_arr[12187] = 8'b00100000;
		color_arr[12188] = 8'b00100000;
		color_arr[12189] = 8'b00100000;
		color_arr[12190] = 8'b00100000;
		color_arr[12191] = 8'b00100000;
		color_arr[12192] = 8'b00100000;
		color_arr[12193] = 8'b00100000;
		color_arr[12194] = 8'b00100000;
		color_arr[12195] = 8'b00100000;
		color_arr[12196] = 8'b00100000;
		color_arr[12197] = 8'b00100000;
		color_arr[12198] = 8'b00100000;
		color_arr[12199] = 8'b00100000;
		color_arr[12200] = 8'b00000000;
		color_arr[12201] = 8'b00000000;
		color_arr[12202] = 8'b00000000;
		color_arr[12203] = 8'b00100000;
		color_arr[12204] = 8'b00100000;
		color_arr[12205] = 8'b00100000;
		color_arr[12206] = 8'b00100000;
		color_arr[12207] = 8'b00100000;
		color_arr[12208] = 8'b00100000;
		color_arr[12209] = 8'b00100000;
		color_arr[12210] = 8'b00100000;
		color_arr[12211] = 8'b00100000;
		color_arr[12212] = 8'b00100000;
		color_arr[12213] = 8'b00100000;
		color_arr[12214] = 8'b00100000;
		color_arr[12215] = 8'b00100000;
		color_arr[12216] = 8'b00100000;
		color_arr[12217] = 8'b00100000;
		color_arr[12218] = 8'b00100000;
		color_arr[12219] = 8'b00100000;
		color_arr[12220] = 8'b00100000;
		color_arr[12221] = 8'b00100000;
		color_arr[12222] = 8'b00000000;
		color_arr[12223] = 8'b00000000;
		color_arr[12224] = 8'b00000000;
		color_arr[12225] = 8'b00000000;
		color_arr[12226] = 8'b00100000;
		color_arr[12227] = 8'b00100000;
		color_arr[12228] = 8'b00100000;
		color_arr[12229] = 8'b00100000;
		color_arr[12230] = 8'b00100000;
		color_arr[12231] = 8'b00100000;
		color_arr[12232] = 8'b00100000;
		color_arr[12233] = 8'b00100000;
		color_arr[12234] = 8'b00100000;
		color_arr[12235] = 8'b00100000;
		color_arr[12236] = 8'b00100000;
		color_arr[12237] = 8'b00100000;
		color_arr[12238] = 8'b00100000;
		color_arr[12239] = 8'b00100000;
		color_arr[12240] = 8'b00001000;
		color_arr[12241] = 8'b00001000;
		color_arr[12242] = 8'b00001000;
		color_arr[12243] = 8'b00001000;
		color_arr[12244] = 8'b00001000;
		color_arr[12245] = 8'b00001000;
		color_arr[12246] = 8'b00001000;
		color_arr[12247] = 8'b00001000;
		color_arr[12248] = 8'b00001000;
		color_arr[12249] = 8'b00001000;
		color_arr[12250] = 8'b00001000;
		color_arr[12251] = 8'b00001000;
		color_arr[12252] = 8'b00001000;
		color_arr[12253] = 8'b00001000;
		color_arr[12254] = 8'b00001000;
		color_arr[12255] = 8'b00001000;
		color_arr[12256] = 8'b00001000;
		color_arr[12257] = 8'b00001000;
		color_arr[12258] = 8'b00001000;
		color_arr[12259] = 8'b00001000;
		color_arr[12260] = 8'b00001000;
		color_arr[12261] = 8'b00001000;
		color_arr[12262] = 8'b00001000;
		color_arr[12263] = 8'b00001000;
		color_arr[12264] = 8'b00001000;
		color_arr[12265] = 8'b00001000;
		color_arr[12266] = 8'b00001000;
		color_arr[12267] = 8'b00001000;
		color_arr[12268] = 8'b00001000;
		color_arr[12269] = 8'b00001000;
		color_arr[12270] = 8'b00001000;
		color_arr[12271] = 8'b00001000;
		color_arr[12272] = 8'b00000000;
		color_arr[12273] = 8'b00000000;
		color_arr[12274] = 8'b00000000;
		color_arr[12275] = 8'b00001000;
		color_arr[12276] = 8'b00001000;
		color_arr[12277] = 8'b00001000;
		color_arr[12278] = 8'b00001000;
		color_arr[12279] = 8'b00000000;
		color_arr[12280] = 8'b00000000;
		color_arr[12281] = 8'b00000000;
		color_arr[12282] = 8'b00001000;
		color_arr[12283] = 8'b00001000;
		color_arr[12284] = 8'b00001000;
		color_arr[12285] = 8'b00010010;
		color_arr[12286] = 8'b00010010;
		color_arr[12287] = 8'b00010010;
		color_arr[12288] = 8'b00010010;
		color_arr[12289] = 8'b00010010;
		color_arr[12290] = 8'b00010010;
		color_arr[12291] = 8'b00010010;
		color_arr[12292] = 8'b00010010;
		color_arr[12293] = 8'b00010010;
		color_arr[12294] = 8'b00010010;
		color_arr[12295] = 8'b00010010;
		color_arr[12296] = 8'b00010010;
		color_arr[12297] = 8'b00010010;
		color_arr[12298] = 8'b00010010;
		color_arr[12299] = 8'b00010010;
		color_arr[12300] = 8'b00010010;
		color_arr[12301] = 8'b00010010;
		color_arr[12302] = 8'b00010010;
		color_arr[12303] = 8'b00010010;
		color_arr[12304] = 8'b00010010;
		color_arr[12305] = 8'b00010010;
		color_arr[12306] = 8'b00100000;
		color_arr[12307] = 8'b00100000;
		color_arr[12308] = 8'b00100000;
		color_arr[12309] = 8'b00100000;
		color_arr[12310] = 8'b00000000;
		color_arr[12311] = 8'b00000000;
		color_arr[12312] = 8'b00100000;
		color_arr[12313] = 8'b00100000;
		color_arr[12314] = 8'b00100000;
		color_arr[12315] = 8'b00100000;
		color_arr[12316] = 8'b00100000;
		color_arr[12317] = 8'b00100000;
		color_arr[12318] = 8'b00100000;
		color_arr[12319] = 8'b00100000;
		color_arr[12320] = 8'b00100000;
		color_arr[12321] = 8'b00100000;
		color_arr[12322] = 8'b00100000;
		color_arr[12323] = 8'b00100000;
		color_arr[12324] = 8'b00100000;
		color_arr[12325] = 8'b00100000;
		color_arr[12326] = 8'b00000000;
		color_arr[12327] = 8'b00000000;
		color_arr[12328] = 8'b00000000;
		color_arr[12329] = 8'b00000000;
		color_arr[12330] = 8'b00100000;
		color_arr[12331] = 8'b00100000;
		color_arr[12332] = 8'b00100000;
		color_arr[12333] = 8'b00100000;
		color_arr[12334] = 8'b00100000;
		color_arr[12335] = 8'b00100000;
		color_arr[12336] = 8'b00100000;
		color_arr[12337] = 8'b00100000;
		color_arr[12338] = 8'b00100000;
		color_arr[12339] = 8'b00100000;
		color_arr[12340] = 8'b00100000;
		color_arr[12341] = 8'b00100000;
		color_arr[12342] = 8'b00100000;
		color_arr[12343] = 8'b00100000;
		color_arr[12344] = 8'b00100000;
		color_arr[12345] = 8'b00100000;
		color_arr[12346] = 8'b00100000;
		color_arr[12347] = 8'b00100000;
		color_arr[12348] = 8'b00100000;
		color_arr[12349] = 8'b00000000;
		color_arr[12350] = 8'b00000000;
		color_arr[12351] = 8'b00000000;
		color_arr[12352] = 8'b00000000;
		color_arr[12353] = 8'b00100000;
		color_arr[12354] = 8'b00100000;
		color_arr[12355] = 8'b00100000;
		color_arr[12356] = 8'b00100000;
		color_arr[12357] = 8'b00100000;
		color_arr[12358] = 8'b00100000;
		color_arr[12359] = 8'b00100000;
		color_arr[12360] = 8'b00100000;
		color_arr[12361] = 8'b00100000;
		color_arr[12362] = 8'b00100000;
		color_arr[12363] = 8'b00100000;
		color_arr[12364] = 8'b00100000;
		color_arr[12365] = 8'b00100000;
		color_arr[12366] = 8'b00100000;
		color_arr[12367] = 8'b00100000;
		color_arr[12368] = 8'b00001000;
		color_arr[12369] = 8'b00001000;
		color_arr[12370] = 8'b00001000;
		color_arr[12371] = 8'b00001000;
		color_arr[12372] = 8'b00001000;
		color_arr[12373] = 8'b00001000;
		color_arr[12374] = 8'b00001000;
		color_arr[12375] = 8'b00001000;
		color_arr[12376] = 8'b00001000;
		color_arr[12377] = 8'b00001000;
		color_arr[12378] = 8'b00001000;
		color_arr[12379] = 8'b00001000;
		color_arr[12380] = 8'b00001000;
		color_arr[12381] = 8'b00001000;
		color_arr[12382] = 8'b00001000;
		color_arr[12383] = 8'b00001000;
		color_arr[12384] = 8'b00001000;
		color_arr[12385] = 8'b00001000;
		color_arr[12386] = 8'b00001000;
		color_arr[12387] = 8'b00001000;
		color_arr[12388] = 8'b00001000;
		color_arr[12389] = 8'b00001000;
		color_arr[12390] = 8'b00001000;
		color_arr[12391] = 8'b00001000;
		color_arr[12392] = 8'b00001000;
		color_arr[12393] = 8'b00001000;
		color_arr[12394] = 8'b00001000;
		color_arr[12395] = 8'b00001000;
		color_arr[12396] = 8'b00001000;
		color_arr[12397] = 8'b00001000;
		color_arr[12398] = 8'b00000000;
		color_arr[12399] = 8'b00000000;
		color_arr[12400] = 8'b00000000;
		color_arr[12401] = 8'b00000000;
		color_arr[12402] = 8'b00001000;
		color_arr[12403] = 8'b00001000;
		color_arr[12404] = 8'b00001000;
		color_arr[12405] = 8'b00001000;
		color_arr[12406] = 8'b00001000;
		color_arr[12407] = 8'b00001000;
		color_arr[12408] = 8'b00000000;
		color_arr[12409] = 8'b00000000;
		color_arr[12410] = 8'b00001000;
		color_arr[12411] = 8'b00001000;
		color_arr[12412] = 8'b00001000;
		color_arr[12413] = 8'b00010010;
		color_arr[12414] = 8'b00010010;
		color_arr[12415] = 8'b00010010;
		color_arr[12416] = 8'b00010010;
		color_arr[12417] = 8'b00010010;
		color_arr[12418] = 8'b00010010;
		color_arr[12419] = 8'b00010010;
		color_arr[12420] = 8'b00010010;
		color_arr[12421] = 8'b00010010;
		color_arr[12422] = 8'b00010010;
		color_arr[12423] = 8'b00010010;
		color_arr[12424] = 8'b00010010;
		color_arr[12425] = 8'b00010010;
		color_arr[12426] = 8'b00010010;
		color_arr[12427] = 8'b00010010;
		color_arr[12428] = 8'b00010010;
		color_arr[12429] = 8'b00010010;
		color_arr[12430] = 8'b00010010;
		color_arr[12431] = 8'b00010010;
		color_arr[12432] = 8'b00010010;
		color_arr[12433] = 8'b00010010;
		color_arr[12434] = 8'b00100000;
		color_arr[12435] = 8'b00100000;
		color_arr[12436] = 8'b00100000;
		color_arr[12437] = 8'b00100000;
		color_arr[12438] = 8'b00000000;
		color_arr[12439] = 8'b00000000;
		color_arr[12440] = 8'b00100000;
		color_arr[12441] = 8'b00100000;
		color_arr[12442] = 8'b00100000;
		color_arr[12443] = 8'b00100000;
		color_arr[12444] = 8'b00100000;
		color_arr[12445] = 8'b00100000;
		color_arr[12446] = 8'b00100000;
		color_arr[12447] = 8'b00100000;
		color_arr[12448] = 8'b00100000;
		color_arr[12449] = 8'b00100000;
		color_arr[12450] = 8'b00100000;
		color_arr[12451] = 8'b00100000;
		color_arr[12452] = 8'b00100000;
		color_arr[12453] = 8'b00000000;
		color_arr[12454] = 8'b00000000;
		color_arr[12455] = 8'b00000000;
		color_arr[12456] = 8'b00000000;
		color_arr[12457] = 8'b00100000;
		color_arr[12458] = 8'b00100000;
		color_arr[12459] = 8'b00100000;
		color_arr[12460] = 8'b00100000;
		color_arr[12461] = 8'b00100000;
		color_arr[12462] = 8'b00100000;
		color_arr[12463] = 8'b00100000;
		color_arr[12464] = 8'b00100000;
		color_arr[12465] = 8'b00100000;
		color_arr[12466] = 8'b00100000;
		color_arr[12467] = 8'b00100000;
		color_arr[12468] = 8'b00100000;
		color_arr[12469] = 8'b00100000;
		color_arr[12470] = 8'b00100000;
		color_arr[12471] = 8'b00100000;
		color_arr[12472] = 8'b00100000;
		color_arr[12473] = 8'b00100000;
		color_arr[12474] = 8'b00100000;
		color_arr[12475] = 8'b00000000;
		color_arr[12476] = 8'b00000000;
		color_arr[12477] = 8'b00000000;
		color_arr[12478] = 8'b00000000;
		color_arr[12479] = 8'b00100000;
		color_arr[12480] = 8'b00100000;
		color_arr[12481] = 8'b00100000;
		color_arr[12482] = 8'b00100000;
		color_arr[12483] = 8'b00100000;
		color_arr[12484] = 8'b00100000;
		color_arr[12485] = 8'b00100000;
		color_arr[12486] = 8'b00100000;
		color_arr[12487] = 8'b00100000;
		color_arr[12488] = 8'b00100000;
		color_arr[12489] = 8'b00100000;
		color_arr[12490] = 8'b00100000;
		color_arr[12491] = 8'b00100000;
		color_arr[12492] = 8'b00100000;
		color_arr[12493] = 8'b00100000;
		color_arr[12494] = 8'b00100000;
		color_arr[12495] = 8'b00100000;
		color_arr[12496] = 8'b00100000;
		color_arr[12497] = 8'b00100000;
		color_arr[12498] = 8'b00100000;
		color_arr[12499] = 8'b00100000;
		color_arr[12500] = 8'b00100000;
		color_arr[12501] = 8'b00100000;
		color_arr[12502] = 8'b00100000;
		color_arr[12503] = 8'b00100000;
		color_arr[12504] = 8'b00100000;
		color_arr[12505] = 8'b00100000;
		color_arr[12506] = 8'b00100000;
		color_arr[12507] = 8'b00100000;
		color_arr[12508] = 8'b00100000;
		color_arr[12509] = 8'b00100000;
		color_arr[12510] = 8'b00100000;
		color_arr[12511] = 8'b00100000;
		color_arr[12512] = 8'b00100000;
		color_arr[12513] = 8'b00100000;
		color_arr[12514] = 8'b00100000;
		color_arr[12515] = 8'b00100000;
		color_arr[12516] = 8'b00100000;
		color_arr[12517] = 8'b00100000;
		color_arr[12518] = 8'b00100000;
		color_arr[12519] = 8'b00100000;
		color_arr[12520] = 8'b00100000;
		color_arr[12521] = 8'b00100000;
		color_arr[12522] = 8'b00100000;
		color_arr[12523] = 8'b00100000;
		color_arr[12524] = 8'b00100000;
		color_arr[12525] = 8'b00000000;
		color_arr[12526] = 8'b00000000;
		color_arr[12527] = 8'b00000000;
		color_arr[12528] = 8'b00000000;
		color_arr[12529] = 8'b00100000;
		color_arr[12530] = 8'b00100000;
		color_arr[12531] = 8'b00100000;
		color_arr[12532] = 8'b00100000;
		color_arr[12533] = 8'b00100000;
		color_arr[12534] = 8'b00100000;
		color_arr[12535] = 8'b00100000;
		color_arr[12536] = 8'b00000000;
		color_arr[12537] = 8'b00000000;
		color_arr[12538] = 8'b00100000;
		color_arr[12539] = 8'b00100000;
		color_arr[12540] = 8'b00100000;
		color_arr[12541] = 8'b00010010;
		color_arr[12542] = 8'b00010010;
		color_arr[12543] = 8'b00010010;
		color_arr[12544] = 8'b00010010;
		color_arr[12545] = 8'b00010010;
		color_arr[12546] = 8'b00010010;
		color_arr[12547] = 8'b00010010;
		color_arr[12548] = 8'b00010010;
		color_arr[12549] = 8'b00010010;
		color_arr[12550] = 8'b00010010;
		color_arr[12551] = 8'b00010010;
		color_arr[12552] = 8'b00010010;
		color_arr[12553] = 8'b00010010;
		color_arr[12554] = 8'b00010010;
		color_arr[12555] = 8'b00010010;
		color_arr[12556] = 8'b00010010;
		color_arr[12557] = 8'b00010010;
		color_arr[12558] = 8'b00010010;
		color_arr[12559] = 8'b00010010;
		color_arr[12560] = 8'b00010010;
		color_arr[12561] = 8'b00010010;
		color_arr[12562] = 8'b00100000;
		color_arr[12563] = 8'b00100000;
		color_arr[12564] = 8'b00100000;
		color_arr[12565] = 8'b00100000;
		color_arr[12566] = 8'b00000000;
		color_arr[12567] = 8'b00000000;
		color_arr[12568] = 8'b00100000;
		color_arr[12569] = 8'b00100000;
		color_arr[12570] = 8'b00100000;
		color_arr[12571] = 8'b00100000;
		color_arr[12572] = 8'b00100000;
		color_arr[12573] = 8'b00100000;
		color_arr[12574] = 8'b00100000;
		color_arr[12575] = 8'b00100000;
		color_arr[12576] = 8'b00100000;
		color_arr[12577] = 8'b00100000;
		color_arr[12578] = 8'b00100000;
		color_arr[12579] = 8'b00000000;
		color_arr[12580] = 8'b00000000;
		color_arr[12581] = 8'b00000000;
		color_arr[12582] = 8'b00000000;
		color_arr[12583] = 8'b00100000;
		color_arr[12584] = 8'b00100000;
		color_arr[12585] = 8'b00100000;
		color_arr[12586] = 8'b00100000;
		color_arr[12587] = 8'b00100000;
		color_arr[12588] = 8'b00100000;
		color_arr[12589] = 8'b00100000;
		color_arr[12590] = 8'b00100000;
		color_arr[12591] = 8'b00100000;
		color_arr[12592] = 8'b00100000;
		color_arr[12593] = 8'b00100000;
		color_arr[12594] = 8'b00100000;
		color_arr[12595] = 8'b00100000;
		color_arr[12596] = 8'b00100000;
		color_arr[12597] = 8'b00100000;
		color_arr[12598] = 8'b00100000;
		color_arr[12599] = 8'b00100000;
		color_arr[12600] = 8'b00100000;
		color_arr[12601] = 8'b00100000;
		color_arr[12602] = 8'b00000000;
		color_arr[12603] = 8'b00000000;
		color_arr[12604] = 8'b00000000;
		color_arr[12605] = 8'b00000000;
		color_arr[12606] = 8'b00100000;
		color_arr[12607] = 8'b00100000;
		color_arr[12608] = 8'b00100000;
		color_arr[12609] = 8'b00100000;
		color_arr[12610] = 8'b00100000;
		color_arr[12611] = 8'b00100000;
		color_arr[12612] = 8'b00100000;
		color_arr[12613] = 8'b00100000;
		color_arr[12614] = 8'b00100000;
		color_arr[12615] = 8'b00100000;
		color_arr[12616] = 8'b00100000;
		color_arr[12617] = 8'b00100000;
		color_arr[12618] = 8'b00100000;
		color_arr[12619] = 8'b00100000;
		color_arr[12620] = 8'b00100000;
		color_arr[12621] = 8'b00100000;
		color_arr[12622] = 8'b00100000;
		color_arr[12623] = 8'b00100000;
		color_arr[12624] = 8'b00100000;
		color_arr[12625] = 8'b00100000;
		color_arr[12626] = 8'b00100000;
		color_arr[12627] = 8'b00100000;
		color_arr[12628] = 8'b00100000;
		color_arr[12629] = 8'b00100000;
		color_arr[12630] = 8'b00100000;
		color_arr[12631] = 8'b00100000;
		color_arr[12632] = 8'b00100000;
		color_arr[12633] = 8'b00100000;
		color_arr[12634] = 8'b00100000;
		color_arr[12635] = 8'b00100000;
		color_arr[12636] = 8'b00100000;
		color_arr[12637] = 8'b00100000;
		color_arr[12638] = 8'b00100000;
		color_arr[12639] = 8'b00100000;
		color_arr[12640] = 8'b00100000;
		color_arr[12641] = 8'b00100000;
		color_arr[12642] = 8'b00100000;
		color_arr[12643] = 8'b00100000;
		color_arr[12644] = 8'b00100000;
		color_arr[12645] = 8'b00100000;
		color_arr[12646] = 8'b00100000;
		color_arr[12647] = 8'b00100000;
		color_arr[12648] = 8'b00100000;
		color_arr[12649] = 8'b00100000;
		color_arr[12650] = 8'b00100000;
		color_arr[12651] = 8'b00100000;
		color_arr[12652] = 8'b00000000;
		color_arr[12653] = 8'b00000000;
		color_arr[12654] = 8'b00000000;
		color_arr[12655] = 8'b00100000;
		color_arr[12656] = 8'b00100000;
		color_arr[12657] = 8'b00100000;
		color_arr[12658] = 8'b00100000;
		color_arr[12659] = 8'b00100000;
		color_arr[12660] = 8'b00100000;
		color_arr[12661] = 8'b00100000;
		color_arr[12662] = 8'b00100000;
		color_arr[12663] = 8'b00100000;
		color_arr[12664] = 8'b00000000;
		color_arr[12665] = 8'b00000000;
		color_arr[12666] = 8'b00100000;
		color_arr[12667] = 8'b00100000;
		color_arr[12668] = 8'b00100000;
		color_arr[12669] = 8'b00010010;
		color_arr[12670] = 8'b00010010;
		color_arr[12671] = 8'b00010010;
		color_arr[12672] = 8'b00010010;
		color_arr[12673] = 8'b00010010;
		color_arr[12674] = 8'b00010010;
		color_arr[12675] = 8'b00010010;
		color_arr[12676] = 8'b00010010;
		color_arr[12677] = 8'b00010010;
		color_arr[12678] = 8'b00010010;
		color_arr[12679] = 8'b00010010;
		color_arr[12680] = 8'b00010010;
		color_arr[12681] = 8'b00010010;
		color_arr[12682] = 8'b00010010;
		color_arr[12683] = 8'b00010010;
		color_arr[12684] = 8'b00010010;
		color_arr[12685] = 8'b00010010;
		color_arr[12686] = 8'b00010010;
		color_arr[12687] = 8'b00010010;
		color_arr[12688] = 8'b00010010;
		color_arr[12689] = 8'b00010010;
		color_arr[12690] = 8'b00100000;
		color_arr[12691] = 8'b00100000;
		color_arr[12692] = 8'b00100000;
		color_arr[12693] = 8'b00100000;
		color_arr[12694] = 8'b00000000;
		color_arr[12695] = 8'b00000000;
		color_arr[12696] = 8'b00100000;
		color_arr[12697] = 8'b00100000;
		color_arr[12698] = 8'b00100000;
		color_arr[12699] = 8'b00100000;
		color_arr[12700] = 8'b00100000;
		color_arr[12701] = 8'b00100000;
		color_arr[12702] = 8'b00100000;
		color_arr[12703] = 8'b00100000;
		color_arr[12704] = 8'b00100000;
		color_arr[12705] = 8'b00000000;
		color_arr[12706] = 8'b00000000;
		color_arr[12707] = 8'b00000000;
		color_arr[12708] = 8'b00000000;
		color_arr[12709] = 8'b00000000;
		color_arr[12710] = 8'b00100000;
		color_arr[12711] = 8'b00100000;
		color_arr[12712] = 8'b00100000;
		color_arr[12713] = 8'b00100000;
		color_arr[12714] = 8'b00100000;
		color_arr[12715] = 8'b00100000;
		color_arr[12716] = 8'b00100000;
		color_arr[12717] = 8'b00100000;
		color_arr[12718] = 8'b00100000;
		color_arr[12719] = 8'b00100000;
		color_arr[12720] = 8'b00100000;
		color_arr[12721] = 8'b00100000;
		color_arr[12722] = 8'b00100000;
		color_arr[12723] = 8'b00100000;
		color_arr[12724] = 8'b00100000;
		color_arr[12725] = 8'b00100000;
		color_arr[12726] = 8'b00100000;
		color_arr[12727] = 8'b00100000;
		color_arr[12728] = 8'b00000000;
		color_arr[12729] = 8'b00000000;
		color_arr[12730] = 8'b00000000;
		color_arr[12731] = 8'b00000000;
		color_arr[12732] = 8'b00000000;
		color_arr[12733] = 8'b00000000;
		color_arr[12734] = 8'b00000000;
		color_arr[12735] = 8'b00000000;
		color_arr[12736] = 8'b00000000;
		color_arr[12737] = 8'b00000000;
		color_arr[12738] = 8'b00000000;
		color_arr[12739] = 8'b00100000;
		color_arr[12740] = 8'b00100000;
		color_arr[12741] = 8'b00100000;
		color_arr[12742] = 8'b00100000;
		color_arr[12743] = 8'b00100000;
		color_arr[12744] = 8'b00100000;
		color_arr[12745] = 8'b00100000;
		color_arr[12746] = 8'b00100000;
		color_arr[12747] = 8'b00100000;
		color_arr[12748] = 8'b00100000;
		color_arr[12749] = 8'b00100000;
		color_arr[12750] = 8'b00100000;
		color_arr[12751] = 8'b00100000;
		color_arr[12752] = 8'b00100000;
		color_arr[12753] = 8'b00100000;
		color_arr[12754] = 8'b00100000;
		color_arr[12755] = 8'b00100000;
		color_arr[12756] = 8'b00100000;
		color_arr[12757] = 8'b00100000;
		color_arr[12758] = 8'b00100000;
		color_arr[12759] = 8'b00100000;
		color_arr[12760] = 8'b00100000;
		color_arr[12761] = 8'b00100000;
		color_arr[12762] = 8'b00100000;
		color_arr[12763] = 8'b00100000;
		color_arr[12764] = 8'b00100000;
		color_arr[12765] = 8'b00100000;
		color_arr[12766] = 8'b00100000;
		color_arr[12767] = 8'b00100000;
		color_arr[12768] = 8'b00100000;
		color_arr[12769] = 8'b00100000;
		color_arr[12770] = 8'b00100000;
		color_arr[12771] = 8'b00100000;
		color_arr[12772] = 8'b00100000;
		color_arr[12773] = 8'b00100000;
		color_arr[12774] = 8'b00100000;
		color_arr[12775] = 8'b00100000;
		color_arr[12776] = 8'b00100000;
		color_arr[12777] = 8'b00100000;
		color_arr[12778] = 8'b00000000;
		color_arr[12779] = 8'b00000000;
		color_arr[12780] = 8'b00000000;
		color_arr[12781] = 8'b00000000;
		color_arr[12782] = 8'b00100000;
		color_arr[12783] = 8'b00100000;
		color_arr[12784] = 8'b00100000;
		color_arr[12785] = 8'b00100000;
		color_arr[12786] = 8'b00100000;
		color_arr[12787] = 8'b00100000;
		color_arr[12788] = 8'b00100000;
		color_arr[12789] = 8'b00100000;
		color_arr[12790] = 8'b00100000;
		color_arr[12791] = 8'b00100000;
		color_arr[12792] = 8'b00000000;
		color_arr[12793] = 8'b00000000;
		color_arr[12794] = 8'b00100000;
		color_arr[12795] = 8'b00100000;
		color_arr[12796] = 8'b00100000;
		color_arr[12797] = 8'b00010010;
		color_arr[12798] = 8'b00010010;
		color_arr[12799] = 8'b00010010;
		color_arr[12800] = 8'b00010010;
		color_arr[12801] = 8'b00010010;
		color_arr[12802] = 8'b00010010;
		color_arr[12803] = 8'b00010010;
		color_arr[12804] = 8'b00010010;
		color_arr[12805] = 8'b00010010;
		color_arr[12806] = 8'b00010010;
		color_arr[12807] = 8'b00010010;
		color_arr[12808] = 8'b00010010;
		color_arr[12809] = 8'b00010010;
		color_arr[12810] = 8'b00010010;
		color_arr[12811] = 8'b00010010;
		color_arr[12812] = 8'b00010010;
		color_arr[12813] = 8'b00010010;
		color_arr[12814] = 8'b00010010;
		color_arr[12815] = 8'b00010010;
		color_arr[12816] = 8'b00010010;
		color_arr[12817] = 8'b00010010;
		color_arr[12818] = 8'b00100000;
		color_arr[12819] = 8'b00100000;
		color_arr[12820] = 8'b00100000;
		color_arr[12821] = 8'b00100000;
		color_arr[12822] = 8'b00000000;
		color_arr[12823] = 8'b00000000;
		color_arr[12824] = 8'b00100000;
		color_arr[12825] = 8'b00100000;
		color_arr[12826] = 8'b00100000;
		color_arr[12827] = 8'b00100000;
		color_arr[12828] = 8'b00100000;
		color_arr[12829] = 8'b00100000;
		color_arr[12830] = 8'b00100000;
		color_arr[12831] = 8'b00000000;
		color_arr[12832] = 8'b00000000;
		color_arr[12833] = 8'b00000000;
		color_arr[12834] = 8'b00000000;
		color_arr[12835] = 8'b00000000;
		color_arr[12836] = 8'b00100000;
		color_arr[12837] = 8'b00100000;
		color_arr[12838] = 8'b00100000;
		color_arr[12839] = 8'b00100000;
		color_arr[12840] = 8'b00100000;
		color_arr[12841] = 8'b00100000;
		color_arr[12842] = 8'b00100000;
		color_arr[12843] = 8'b00100000;
		color_arr[12844] = 8'b00100000;
		color_arr[12845] = 8'b00100000;
		color_arr[12846] = 8'b00100000;
		color_arr[12847] = 8'b00100000;
		color_arr[12848] = 8'b00100000;
		color_arr[12849] = 8'b00100000;
		color_arr[12850] = 8'b00100000;
		color_arr[12851] = 8'b00100000;
		color_arr[12852] = 8'b00100000;
		color_arr[12853] = 8'b00000000;
		color_arr[12854] = 8'b00000000;
		color_arr[12855] = 8'b00000000;
		color_arr[12856] = 8'b00000000;
		color_arr[12857] = 8'b00000000;
		color_arr[12858] = 8'b00000000;
		color_arr[12859] = 8'b00000000;
		color_arr[12860] = 8'b00000000;
		color_arr[12861] = 8'b00000000;
		color_arr[12862] = 8'b00000000;
		color_arr[12863] = 8'b00000000;
		color_arr[12864] = 8'b00000000;
		color_arr[12865] = 8'b00000000;
		color_arr[12866] = 8'b00000000;
		color_arr[12867] = 8'b00000000;
		color_arr[12868] = 8'b00000000;
		color_arr[12869] = 8'b00000000;
		color_arr[12870] = 8'b00000000;
		color_arr[12871] = 8'b00100000;
		color_arr[12872] = 8'b00100000;
		color_arr[12873] = 8'b00100000;
		color_arr[12874] = 8'b00100000;
		color_arr[12875] = 8'b00100000;
		color_arr[12876] = 8'b00100000;
		color_arr[12877] = 8'b00100000;
		color_arr[12878] = 8'b00100000;
		color_arr[12879] = 8'b00100000;
		color_arr[12880] = 8'b00100000;
		color_arr[12881] = 8'b00100000;
		color_arr[12882] = 8'b00100000;
		color_arr[12883] = 8'b00100000;
		color_arr[12884] = 8'b00100000;
		color_arr[12885] = 8'b00100000;
		color_arr[12886] = 8'b00100000;
		color_arr[12887] = 8'b00100000;
		color_arr[12888] = 8'b00100000;
		color_arr[12889] = 8'b00100000;
		color_arr[12890] = 8'b00100000;
		color_arr[12891] = 8'b00100000;
		color_arr[12892] = 8'b00100000;
		color_arr[12893] = 8'b00100000;
		color_arr[12894] = 8'b00100000;
		color_arr[12895] = 8'b00100000;
		color_arr[12896] = 8'b00100000;
		color_arr[12897] = 8'b00100000;
		color_arr[12898] = 8'b00100000;
		color_arr[12899] = 8'b00100000;
		color_arr[12900] = 8'b00100000;
		color_arr[12901] = 8'b00100000;
		color_arr[12902] = 8'b00100000;
		color_arr[12903] = 8'b00100000;
		color_arr[12904] = 8'b00100000;
		color_arr[12905] = 8'b00000000;
		color_arr[12906] = 8'b00000000;
		color_arr[12907] = 8'b00000000;
		color_arr[12908] = 8'b00000000;
		color_arr[12909] = 8'b00100000;
		color_arr[12910] = 8'b00100000;
		color_arr[12911] = 8'b00100000;
		color_arr[12912] = 8'b00100000;
		color_arr[12913] = 8'b00100000;
		color_arr[12914] = 8'b00100000;
		color_arr[12915] = 8'b00100000;
		color_arr[12916] = 8'b00100000;
		color_arr[12917] = 8'b00100000;
		color_arr[12918] = 8'b00100000;
		color_arr[12919] = 8'b00100000;
		color_arr[12920] = 8'b00000000;
		color_arr[12921] = 8'b00000000;
		color_arr[12922] = 8'b00100000;
		color_arr[12923] = 8'b00100000;
		color_arr[12924] = 8'b00100000;
		color_arr[12925] = 8'b00010010;
		color_arr[12926] = 8'b00010010;
		color_arr[12927] = 8'b00010010;
		color_arr[12928] = 8'b00010010;
		color_arr[12929] = 8'b00010010;
		color_arr[12930] = 8'b00010010;
		color_arr[12931] = 8'b00010010;
		color_arr[12932] = 8'b00010010;
		color_arr[12933] = 8'b00010010;
		color_arr[12934] = 8'b00010010;
		color_arr[12935] = 8'b00010010;
		color_arr[12936] = 8'b00010010;
		color_arr[12937] = 8'b00010010;
		color_arr[12938] = 8'b00010010;
		color_arr[12939] = 8'b00010010;
		color_arr[12940] = 8'b00010010;
		color_arr[12941] = 8'b00010010;
		color_arr[12942] = 8'b00010010;
		color_arr[12943] = 8'b00010010;
		color_arr[12944] = 8'b00010010;
		color_arr[12945] = 8'b00010010;
		color_arr[12946] = 8'b00100000;
		color_arr[12947] = 8'b00100000;
		color_arr[12948] = 8'b00100000;
		color_arr[12949] = 8'b00100000;
		color_arr[12950] = 8'b00000000;
		color_arr[12951] = 8'b00000000;
		color_arr[12952] = 8'b00100000;
		color_arr[12953] = 8'b00100000;
		color_arr[12954] = 8'b00100000;
		color_arr[12955] = 8'b00100000;
		color_arr[12956] = 8'b00000000;
		color_arr[12957] = 8'b00000000;
		color_arr[12958] = 8'b00000000;
		color_arr[12959] = 8'b00000000;
		color_arr[12960] = 8'b00000000;
		color_arr[12961] = 8'b00000000;
		color_arr[12962] = 8'b00100000;
		color_arr[12963] = 8'b00100000;
		color_arr[12964] = 8'b00100000;
		color_arr[12965] = 8'b00100000;
		color_arr[12966] = 8'b00100000;
		color_arr[12967] = 8'b00100000;
		color_arr[12968] = 8'b00100000;
		color_arr[12969] = 8'b00100000;
		color_arr[12970] = 8'b00100000;
		color_arr[12971] = 8'b00100000;
		color_arr[12972] = 8'b00100000;
		color_arr[12973] = 8'b00100000;
		color_arr[12974] = 8'b00100000;
		color_arr[12975] = 8'b00100000;
		color_arr[12976] = 8'b00100000;
		color_arr[12977] = 8'b00100000;
		color_arr[12978] = 8'b00100000;
		color_arr[12979] = 8'b00000000;
		color_arr[12980] = 8'b00000000;
		color_arr[12981] = 8'b00000000;
		color_arr[12982] = 8'b00000000;
		color_arr[12983] = 8'b00000000;
		color_arr[12984] = 8'b00000000;
		color_arr[12985] = 8'b00000000;
		color_arr[12986] = 8'b00000000;
		color_arr[12987] = 8'b00100000;
		color_arr[12988] = 8'b00100000;
		color_arr[12989] = 8'b00100000;
		color_arr[12990] = 8'b00100000;
		color_arr[12991] = 8'b00100000;
		color_arr[12992] = 8'b00100000;
		color_arr[12993] = 8'b00100000;
		color_arr[12994] = 8'b00000000;
		color_arr[12995] = 8'b00000000;
		color_arr[12996] = 8'b00000000;
		color_arr[12997] = 8'b00000000;
		color_arr[12998] = 8'b00000000;
		color_arr[12999] = 8'b00000000;
		color_arr[13000] = 8'b00100000;
		color_arr[13001] = 8'b00100000;
		color_arr[13002] = 8'b00100000;
		color_arr[13003] = 8'b00100000;
		color_arr[13004] = 8'b00100000;
		color_arr[13005] = 8'b00100000;
		color_arr[13006] = 8'b00100000;
		color_arr[13007] = 8'b00100000;
		color_arr[13008] = 8'b00100000;
		color_arr[13009] = 8'b00100000;
		color_arr[13010] = 8'b00100000;
		color_arr[13011] = 8'b00100000;
		color_arr[13012] = 8'b00100000;
		color_arr[13013] = 8'b00100000;
		color_arr[13014] = 8'b00100000;
		color_arr[13015] = 8'b00100000;
		color_arr[13016] = 8'b00100000;
		color_arr[13017] = 8'b00100000;
		color_arr[13018] = 8'b00100000;
		color_arr[13019] = 8'b00100000;
		color_arr[13020] = 8'b00100000;
		color_arr[13021] = 8'b00100000;
		color_arr[13022] = 8'b00100000;
		color_arr[13023] = 8'b00100000;
		color_arr[13024] = 8'b00100000;
		color_arr[13025] = 8'b00100000;
		color_arr[13026] = 8'b00100000;
		color_arr[13027] = 8'b00100000;
		color_arr[13028] = 8'b00100000;
		color_arr[13029] = 8'b00100000;
		color_arr[13030] = 8'b00100000;
		color_arr[13031] = 8'b00100000;
		color_arr[13032] = 8'b00000000;
		color_arr[13033] = 8'b00000000;
		color_arr[13034] = 8'b00000000;
		color_arr[13035] = 8'b00100000;
		color_arr[13036] = 8'b00100000;
		color_arr[13037] = 8'b00100000;
		color_arr[13038] = 8'b00100000;
		color_arr[13039] = 8'b00100000;
		color_arr[13040] = 8'b00100000;
		color_arr[13041] = 8'b00100000;
		color_arr[13042] = 8'b00100000;
		color_arr[13043] = 8'b00100000;
		color_arr[13044] = 8'b00100000;
		color_arr[13045] = 8'b00100000;
		color_arr[13046] = 8'b00100000;
		color_arr[13047] = 8'b00100000;
		color_arr[13048] = 8'b00000000;
		color_arr[13049] = 8'b00000000;
		color_arr[13050] = 8'b00100000;
		color_arr[13051] = 8'b00100000;
		color_arr[13052] = 8'b00100000;
		color_arr[13053] = 8'b00010010;
		color_arr[13054] = 8'b00010010;
		color_arr[13055] = 8'b00010010;
		color_arr[13056] = 8'b00010010;
		color_arr[13057] = 8'b00010010;
		color_arr[13058] = 8'b00010010;
		color_arr[13059] = 8'b00010010;
		color_arr[13060] = 8'b00010010;
		color_arr[13061] = 8'b00010010;
		color_arr[13062] = 8'b00010010;
		color_arr[13063] = 8'b00010010;
		color_arr[13064] = 8'b00010010;
		color_arr[13065] = 8'b00010010;
		color_arr[13066] = 8'b00010010;
		color_arr[13067] = 8'b00010010;
		color_arr[13068] = 8'b00010010;
		color_arr[13069] = 8'b00010010;
		color_arr[13070] = 8'b00010010;
		color_arr[13071] = 8'b00010010;
		color_arr[13072] = 8'b00010010;
		color_arr[13073] = 8'b00010010;
		color_arr[13074] = 8'b00100000;
		color_arr[13075] = 8'b00100000;
		color_arr[13076] = 8'b00100000;
		color_arr[13077] = 8'b00100000;
		color_arr[13078] = 8'b00000000;
		color_arr[13079] = 8'b00000000;
		color_arr[13080] = 8'b00100000;
		color_arr[13081] = 8'b00100000;
		color_arr[13082] = 8'b00000000;
		color_arr[13083] = 8'b00000000;
		color_arr[13084] = 8'b00000000;
		color_arr[13085] = 8'b00000000;
		color_arr[13086] = 8'b00000000;
		color_arr[13087] = 8'b00000000;
		color_arr[13088] = 8'b00100000;
		color_arr[13089] = 8'b00100000;
		color_arr[13090] = 8'b00100000;
		color_arr[13091] = 8'b00100000;
		color_arr[13092] = 8'b00100000;
		color_arr[13093] = 8'b00100000;
		color_arr[13094] = 8'b00100000;
		color_arr[13095] = 8'b00100000;
		color_arr[13096] = 8'b00100000;
		color_arr[13097] = 8'b00100000;
		color_arr[13098] = 8'b00100000;
		color_arr[13099] = 8'b00100000;
		color_arr[13100] = 8'b00100000;
		color_arr[13101] = 8'b00100000;
		color_arr[13102] = 8'b00100000;
		color_arr[13103] = 8'b00100000;
		color_arr[13104] = 8'b00100000;
		color_arr[13105] = 8'b00000000;
		color_arr[13106] = 8'b00000000;
		color_arr[13107] = 8'b00000000;
		color_arr[13108] = 8'b00000000;
		color_arr[13109] = 8'b00000000;
		color_arr[13110] = 8'b00000000;
		color_arr[13111] = 8'b00000000;
		color_arr[13112] = 8'b00100000;
		color_arr[13113] = 8'b00100000;
		color_arr[13114] = 8'b00100000;
		color_arr[13115] = 8'b00100000;
		color_arr[13116] = 8'b00100000;
		color_arr[13117] = 8'b00100000;
		color_arr[13118] = 8'b00100000;
		color_arr[13119] = 8'b00100000;
		color_arr[13120] = 8'b00100000;
		color_arr[13121] = 8'b00100000;
		color_arr[13122] = 8'b00100000;
		color_arr[13123] = 8'b00100000;
		color_arr[13124] = 8'b00100000;
		color_arr[13125] = 8'b00100000;
		color_arr[13126] = 8'b00000000;
		color_arr[13127] = 8'b00000000;
		color_arr[13128] = 8'b00000000;
		color_arr[13129] = 8'b00000000;
		color_arr[13130] = 8'b00100000;
		color_arr[13131] = 8'b00100000;
		color_arr[13132] = 8'b00100000;
		color_arr[13133] = 8'b00100000;
		color_arr[13134] = 8'b00100000;
		color_arr[13135] = 8'b00100000;
		color_arr[13136] = 8'b00100000;
		color_arr[13137] = 8'b00100000;
		color_arr[13138] = 8'b00100000;
		color_arr[13139] = 8'b00100000;
		color_arr[13140] = 8'b00100000;
		color_arr[13141] = 8'b00100000;
		color_arr[13142] = 8'b00100000;
		color_arr[13143] = 8'b00100000;
		color_arr[13144] = 8'b00100000;
		color_arr[13145] = 8'b00100000;
		color_arr[13146] = 8'b00100000;
		color_arr[13147] = 8'b00100000;
		color_arr[13148] = 8'b00100000;
		color_arr[13149] = 8'b00100000;
		color_arr[13150] = 8'b00100000;
		color_arr[13151] = 8'b00100000;
		color_arr[13152] = 8'b00100000;
		color_arr[13153] = 8'b00100000;
		color_arr[13154] = 8'b00100000;
		color_arr[13155] = 8'b00100000;
		color_arr[13156] = 8'b00100000;
		color_arr[13157] = 8'b00100000;
		color_arr[13158] = 8'b00000000;
		color_arr[13159] = 8'b00000000;
		color_arr[13160] = 8'b00000000;
		color_arr[13161] = 8'b00000000;
		color_arr[13162] = 8'b00100000;
		color_arr[13163] = 8'b00100000;
		color_arr[13164] = 8'b00100000;
		color_arr[13165] = 8'b00100000;
		color_arr[13166] = 8'b00100000;
		color_arr[13167] = 8'b00100000;
		color_arr[13168] = 8'b00100000;
		color_arr[13169] = 8'b00100000;
		color_arr[13170] = 8'b00100000;
		color_arr[13171] = 8'b00100000;
		color_arr[13172] = 8'b00100000;
		color_arr[13173] = 8'b00100000;
		color_arr[13174] = 8'b00100000;
		color_arr[13175] = 8'b00100000;
		color_arr[13176] = 8'b00000000;
		color_arr[13177] = 8'b00000000;
		color_arr[13178] = 8'b00100000;
		color_arr[13179] = 8'b00100000;
		color_arr[13180] = 8'b00100000;
		color_arr[13181] = 8'b00010010;
		color_arr[13182] = 8'b00010010;
		color_arr[13183] = 8'b00010010;
		color_arr[13184] = 8'b00010010;
		color_arr[13185] = 8'b00010010;
		color_arr[13186] = 8'b00010010;
		color_arr[13187] = 8'b00010010;
		color_arr[13188] = 8'b00010010;
		color_arr[13189] = 8'b00010010;
		color_arr[13190] = 8'b00010010;
		color_arr[13191] = 8'b00010010;
		color_arr[13192] = 8'b00010010;
		color_arr[13193] = 8'b00010010;
		color_arr[13194] = 8'b00010010;
		color_arr[13195] = 8'b00010010;
		color_arr[13196] = 8'b00010010;
		color_arr[13197] = 8'b00010010;
		color_arr[13198] = 8'b00010010;
		color_arr[13199] = 8'b00010010;
		color_arr[13200] = 8'b00010010;
		color_arr[13201] = 8'b00010010;
		color_arr[13202] = 8'b00100000;
		color_arr[13203] = 8'b00100000;
		color_arr[13204] = 8'b00100000;
		color_arr[13205] = 8'b00100000;
		color_arr[13206] = 8'b00000000;
		color_arr[13207] = 8'b00000000;
		color_arr[13208] = 8'b00000000;
		color_arr[13209] = 8'b00000000;
		color_arr[13210] = 8'b00000000;
		color_arr[13211] = 8'b00000000;
		color_arr[13212] = 8'b00000000;
		color_arr[13213] = 8'b00100000;
		color_arr[13214] = 8'b00100000;
		color_arr[13215] = 8'b00100000;
		color_arr[13216] = 8'b00100000;
		color_arr[13217] = 8'b00100000;
		color_arr[13218] = 8'b00100000;
		color_arr[13219] = 8'b00100000;
		color_arr[13220] = 8'b00100000;
		color_arr[13221] = 8'b00100000;
		color_arr[13222] = 8'b00100000;
		color_arr[13223] = 8'b00100000;
		color_arr[13224] = 8'b00100000;
		color_arr[13225] = 8'b00100000;
		color_arr[13226] = 8'b00100000;
		color_arr[13227] = 8'b00100000;
		color_arr[13228] = 8'b00100000;
		color_arr[13229] = 8'b00100000;
		color_arr[13230] = 8'b00100000;
		color_arr[13231] = 8'b00000000;
		color_arr[13232] = 8'b00000000;
		color_arr[13233] = 8'b00000000;
		color_arr[13234] = 8'b00000000;
		color_arr[13235] = 8'b00000000;
		color_arr[13236] = 8'b00000000;
		color_arr[13237] = 8'b00000000;
		color_arr[13238] = 8'b00100000;
		color_arr[13239] = 8'b00100000;
		color_arr[13240] = 8'b00100000;
		color_arr[13241] = 8'b00100000;
		color_arr[13242] = 8'b00100000;
		color_arr[13243] = 8'b00100000;
		color_arr[13244] = 8'b00100000;
		color_arr[13245] = 8'b00100000;
		color_arr[13246] = 8'b00100000;
		color_arr[13247] = 8'b00100000;
		color_arr[13248] = 8'b00100000;
		color_arr[13249] = 8'b00100000;
		color_arr[13250] = 8'b00100000;
		color_arr[13251] = 8'b00100000;
		color_arr[13252] = 8'b00100000;
		color_arr[13253] = 8'b00100000;
		color_arr[13254] = 8'b00100000;
		color_arr[13255] = 8'b00000000;
		color_arr[13256] = 8'b00000000;
		color_arr[13257] = 8'b00000000;
		color_arr[13258] = 8'b00000000;
		color_arr[13259] = 8'b00100000;
		color_arr[13260] = 8'b00100000;
		color_arr[13261] = 8'b00100000;
		color_arr[13262] = 8'b00100000;
		color_arr[13263] = 8'b00100000;
		color_arr[13264] = 8'b00100000;
		color_arr[13265] = 8'b00100000;
		color_arr[13266] = 8'b00100000;
		color_arr[13267] = 8'b00100000;
		color_arr[13268] = 8'b00100000;
		color_arr[13269] = 8'b00100000;
		color_arr[13270] = 8'b00100000;
		color_arr[13271] = 8'b00100000;
		color_arr[13272] = 8'b00100000;
		color_arr[13273] = 8'b00100000;
		color_arr[13274] = 8'b00100000;
		color_arr[13275] = 8'b00100000;
		color_arr[13276] = 8'b00100000;
		color_arr[13277] = 8'b00100000;
		color_arr[13278] = 8'b00100000;
		color_arr[13279] = 8'b00100000;
		color_arr[13280] = 8'b00100000;
		color_arr[13281] = 8'b00100000;
		color_arr[13282] = 8'b00100000;
		color_arr[13283] = 8'b00100000;
		color_arr[13284] = 8'b00000000;
		color_arr[13285] = 8'b00000000;
		color_arr[13286] = 8'b00000000;
		color_arr[13287] = 8'b00000000;
		color_arr[13288] = 8'b00000000;
		color_arr[13289] = 8'b00100000;
		color_arr[13290] = 8'b00100000;
		color_arr[13291] = 8'b00100000;
		color_arr[13292] = 8'b00100000;
		color_arr[13293] = 8'b00100000;
		color_arr[13294] = 8'b00100000;
		color_arr[13295] = 8'b00100000;
		color_arr[13296] = 8'b00100000;
		color_arr[13297] = 8'b00100000;
		color_arr[13298] = 8'b00100000;
		color_arr[13299] = 8'b00100000;
		color_arr[13300] = 8'b00100000;
		color_arr[13301] = 8'b00100000;
		color_arr[13302] = 8'b00100000;
		color_arr[13303] = 8'b00100000;
		color_arr[13304] = 8'b00000000;
		color_arr[13305] = 8'b00000000;
		color_arr[13306] = 8'b00100000;
		color_arr[13307] = 8'b00100000;
		color_arr[13308] = 8'b00100000;
		color_arr[13309] = 8'b00010010;
		color_arr[13310] = 8'b00010010;
		color_arr[13311] = 8'b00010010;
		color_arr[13312] = 8'b00010010;
		color_arr[13313] = 8'b00010010;
		color_arr[13314] = 8'b00010010;
		color_arr[13315] = 8'b00010010;
		color_arr[13316] = 8'b00010010;
		color_arr[13317] = 8'b00010010;
		color_arr[13318] = 8'b00010010;
		color_arr[13319] = 8'b00010010;
		color_arr[13320] = 8'b00010010;
		color_arr[13321] = 8'b00010010;
		color_arr[13322] = 8'b00010010;
		color_arr[13323] = 8'b00010010;
		color_arr[13324] = 8'b00010010;
		color_arr[13325] = 8'b00010010;
		color_arr[13326] = 8'b00010010;
		color_arr[13327] = 8'b00010010;
		color_arr[13328] = 8'b00010010;
		color_arr[13329] = 8'b00010010;
		color_arr[13330] = 8'b00100000;
		color_arr[13331] = 8'b00100000;
		color_arr[13332] = 8'b00100000;
		color_arr[13333] = 8'b00100000;
		color_arr[13334] = 8'b00100000;
		color_arr[13335] = 8'b00000000;
		color_arr[13336] = 8'b00000000;
		color_arr[13337] = 8'b00000000;
		color_arr[13338] = 8'b00000000;
		color_arr[13339] = 8'b00100000;
		color_arr[13340] = 8'b00100000;
		color_arr[13341] = 8'b00100000;
		color_arr[13342] = 8'b00100000;
		color_arr[13343] = 8'b00100000;
		color_arr[13344] = 8'b00100000;
		color_arr[13345] = 8'b00100000;
		color_arr[13346] = 8'b00100000;
		color_arr[13347] = 8'b00100000;
		color_arr[13348] = 8'b00100000;
		color_arr[13349] = 8'b00100000;
		color_arr[13350] = 8'b00100000;
		color_arr[13351] = 8'b00100000;
		color_arr[13352] = 8'b00100000;
		color_arr[13353] = 8'b00100000;
		color_arr[13354] = 8'b00100000;
		color_arr[13355] = 8'b00100000;
		color_arr[13356] = 8'b00100000;
		color_arr[13357] = 8'b00100000;
		color_arr[13358] = 8'b00000000;
		color_arr[13359] = 8'b00000000;
		color_arr[13360] = 8'b00000000;
		color_arr[13361] = 8'b00000000;
		color_arr[13362] = 8'b00000000;
		color_arr[13363] = 8'b00000000;
		color_arr[13364] = 8'b00000000;
		color_arr[13365] = 8'b00100000;
		color_arr[13366] = 8'b00100000;
		color_arr[13367] = 8'b00100000;
		color_arr[13368] = 8'b00100000;
		color_arr[13369] = 8'b00100000;
		color_arr[13370] = 8'b00100000;
		color_arr[13371] = 8'b00100000;
		color_arr[13372] = 8'b00100000;
		color_arr[13373] = 8'b00100000;
		color_arr[13374] = 8'b00100000;
		color_arr[13375] = 8'b00100000;
		color_arr[13376] = 8'b00100000;
		color_arr[13377] = 8'b00100000;
		color_arr[13378] = 8'b00100000;
		color_arr[13379] = 8'b00100000;
		color_arr[13380] = 8'b00100000;
		color_arr[13381] = 8'b00100000;
		color_arr[13382] = 8'b00100000;
		color_arr[13383] = 8'b00100000;
		color_arr[13384] = 8'b00100000;
		color_arr[13385] = 8'b00000000;
		color_arr[13386] = 8'b00000000;
		color_arr[13387] = 8'b00000000;
		color_arr[13388] = 8'b00000000;
		color_arr[13389] = 8'b00100000;
		color_arr[13390] = 8'b00100000;
		color_arr[13391] = 8'b00100000;
		color_arr[13392] = 8'b00100000;
		color_arr[13393] = 8'b00100000;
		color_arr[13394] = 8'b00100000;
		color_arr[13395] = 8'b00100000;
		color_arr[13396] = 8'b00100000;
		color_arr[13397] = 8'b00100000;
		color_arr[13398] = 8'b00100000;
		color_arr[13399] = 8'b00100000;
		color_arr[13400] = 8'b00100000;
		color_arr[13401] = 8'b00100000;
		color_arr[13402] = 8'b00100000;
		color_arr[13403] = 8'b00100000;
		color_arr[13404] = 8'b00100000;
		color_arr[13405] = 8'b00100000;
		color_arr[13406] = 8'b00100000;
		color_arr[13407] = 8'b00100000;
		color_arr[13408] = 8'b00100000;
		color_arr[13409] = 8'b00100000;
		color_arr[13410] = 8'b00000000;
		color_arr[13411] = 8'b00000000;
		color_arr[13412] = 8'b00000000;
		color_arr[13413] = 8'b00000000;
		color_arr[13414] = 8'b00000000;
		color_arr[13415] = 8'b00100000;
		color_arr[13416] = 8'b00100000;
		color_arr[13417] = 8'b00100000;
		color_arr[13418] = 8'b00100000;
		color_arr[13419] = 8'b00100000;
		color_arr[13420] = 8'b00100000;
		color_arr[13421] = 8'b00100000;
		color_arr[13422] = 8'b00100000;
		color_arr[13423] = 8'b00100000;
		color_arr[13424] = 8'b00100000;
		color_arr[13425] = 8'b00100000;
		color_arr[13426] = 8'b00100000;
		color_arr[13427] = 8'b00100000;
		color_arr[13428] = 8'b00100000;
		color_arr[13429] = 8'b00100000;
		color_arr[13430] = 8'b00100000;
		color_arr[13431] = 8'b00100000;
		color_arr[13432] = 8'b00000000;
		color_arr[13433] = 8'b00000000;
		color_arr[13434] = 8'b00100000;
		color_arr[13435] = 8'b00100000;
		color_arr[13436] = 8'b00100000;
		color_arr[13437] = 8'b00010010;
		color_arr[13438] = 8'b00010010;
		color_arr[13439] = 8'b00010010;
		color_arr[13440] = 8'b00010010;
		color_arr[13441] = 8'b00010010;
		color_arr[13442] = 8'b00010010;
		color_arr[13443] = 8'b00010010;
		color_arr[13444] = 8'b00010010;
		color_arr[13445] = 8'b00010010;
		color_arr[13446] = 8'b00010010;
		color_arr[13447] = 8'b00010010;
		color_arr[13448] = 8'b00010010;
		color_arr[13449] = 8'b00010010;
		color_arr[13450] = 8'b00010010;
		color_arr[13451] = 8'b00010010;
		color_arr[13452] = 8'b00010010;
		color_arr[13453] = 8'b00010010;
		color_arr[13454] = 8'b00010010;
		color_arr[13455] = 8'b00010010;
		color_arr[13456] = 8'b00010010;
		color_arr[13457] = 8'b00010010;
		color_arr[13458] = 8'b00100000;
		color_arr[13459] = 8'b00100000;
		color_arr[13460] = 8'b00100000;
		color_arr[13461] = 8'b00100000;
		color_arr[13462] = 8'b00100000;
		color_arr[13463] = 8'b00100000;
		color_arr[13464] = 8'b00100000;
		color_arr[13465] = 8'b00100000;
		color_arr[13466] = 8'b00100000;
		color_arr[13467] = 8'b00100000;
		color_arr[13468] = 8'b00100000;
		color_arr[13469] = 8'b00100000;
		color_arr[13470] = 8'b00100000;
		color_arr[13471] = 8'b00100000;
		color_arr[13472] = 8'b00100000;
		color_arr[13473] = 8'b00100000;
		color_arr[13474] = 8'b00100000;
		color_arr[13475] = 8'b00100000;
		color_arr[13476] = 8'b00100000;
		color_arr[13477] = 8'b00100000;
		color_arr[13478] = 8'b00100000;
		color_arr[13479] = 8'b00100000;
		color_arr[13480] = 8'b00100000;
		color_arr[13481] = 8'b00100000;
		color_arr[13482] = 8'b00100000;
		color_arr[13483] = 8'b00100000;
		color_arr[13484] = 8'b00100000;
		color_arr[13485] = 8'b00000000;
		color_arr[13486] = 8'b00000000;
		color_arr[13487] = 8'b00000000;
		color_arr[13488] = 8'b00000000;
		color_arr[13489] = 8'b00000000;
		color_arr[13490] = 8'b00000000;
		color_arr[13491] = 8'b00000000;
		color_arr[13492] = 8'b00100000;
		color_arr[13493] = 8'b00100000;
		color_arr[13494] = 8'b00100000;
		color_arr[13495] = 8'b00100000;
		color_arr[13496] = 8'b00100000;
		color_arr[13497] = 8'b00100000;
		color_arr[13498] = 8'b00100000;
		color_arr[13499] = 8'b00100000;
		color_arr[13500] = 8'b00100000;
		color_arr[13501] = 8'b00100000;
		color_arr[13502] = 8'b00100000;
		color_arr[13503] = 8'b00100000;
		color_arr[13504] = 8'b00100000;
		color_arr[13505] = 8'b00100000;
		color_arr[13506] = 8'b00100000;
		color_arr[13507] = 8'b00100000;
		color_arr[13508] = 8'b00100000;
		color_arr[13509] = 8'b00100000;
		color_arr[13510] = 8'b00100000;
		color_arr[13511] = 8'b00100000;
		color_arr[13512] = 8'b00100000;
		color_arr[13513] = 8'b00100000;
		color_arr[13514] = 8'b00000000;
		color_arr[13515] = 8'b00000000;
		color_arr[13516] = 8'b00000000;
		color_arr[13517] = 8'b00000000;
		color_arr[13518] = 8'b00100000;
		color_arr[13519] = 8'b00100000;
		color_arr[13520] = 8'b00100000;
		color_arr[13521] = 8'b00100000;
		color_arr[13522] = 8'b00100000;
		color_arr[13523] = 8'b00100000;
		color_arr[13524] = 8'b00100000;
		color_arr[13525] = 8'b00100000;
		color_arr[13526] = 8'b00100000;
		color_arr[13527] = 8'b00100000;
		color_arr[13528] = 8'b00100000;
		color_arr[13529] = 8'b00100000;
		color_arr[13530] = 8'b00100000;
		color_arr[13531] = 8'b00100000;
		color_arr[13532] = 8'b00100000;
		color_arr[13533] = 8'b00100000;
		color_arr[13534] = 8'b00100000;
		color_arr[13535] = 8'b00100000;
		color_arr[13536] = 8'b00000000;
		color_arr[13537] = 8'b00000000;
		color_arr[13538] = 8'b00000000;
		color_arr[13539] = 8'b00000000;
		color_arr[13540] = 8'b00000000;
		color_arr[13541] = 8'b00100000;
		color_arr[13542] = 8'b00100000;
		color_arr[13543] = 8'b00100000;
		color_arr[13544] = 8'b00100000;
		color_arr[13545] = 8'b00100000;
		color_arr[13546] = 8'b00100000;
		color_arr[13547] = 8'b00100000;
		color_arr[13548] = 8'b00100000;
		color_arr[13549] = 8'b00100000;
		color_arr[13550] = 8'b00100000;
		color_arr[13551] = 8'b00100000;
		color_arr[13552] = 8'b00100000;
		color_arr[13553] = 8'b00100000;
		color_arr[13554] = 8'b00100000;
		color_arr[13555] = 8'b00100000;
		color_arr[13556] = 8'b00100000;
		color_arr[13557] = 8'b00100000;
		color_arr[13558] = 8'b00100000;
		color_arr[13559] = 8'b00100000;
		color_arr[13560] = 8'b00000000;
		color_arr[13561] = 8'b00000000;
		color_arr[13562] = 8'b00100000;
		color_arr[13563] = 8'b00100000;
		color_arr[13564] = 8'b00100000;
		color_arr[13565] = 8'b00010010;
		color_arr[13566] = 8'b00010010;
		color_arr[13567] = 8'b00010010;
		color_arr[13568] = 8'b00010010;
		color_arr[13569] = 8'b00010010;
		color_arr[13570] = 8'b00010010;
		color_arr[13571] = 8'b00010010;
		color_arr[13572] = 8'b00010010;
		color_arr[13573] = 8'b00010010;
		color_arr[13574] = 8'b00010010;
		color_arr[13575] = 8'b00010010;
		color_arr[13576] = 8'b00010010;
		color_arr[13577] = 8'b00010010;
		color_arr[13578] = 8'b00010010;
		color_arr[13579] = 8'b00010010;
		color_arr[13580] = 8'b00010010;
		color_arr[13581] = 8'b00010010;
		color_arr[13582] = 8'b00010010;
		color_arr[13583] = 8'b00010010;
		color_arr[13584] = 8'b00010010;
		color_arr[13585] = 8'b00010010;
		color_arr[13586] = 8'b00100000;
		color_arr[13587] = 8'b00100000;
		color_arr[13588] = 8'b00100000;
		color_arr[13589] = 8'b00100000;
		color_arr[13590] = 8'b00100000;
		color_arr[13591] = 8'b00100000;
		color_arr[13592] = 8'b00100000;
		color_arr[13593] = 8'b00100000;
		color_arr[13594] = 8'b00100000;
		color_arr[13595] = 8'b00100000;
		color_arr[13596] = 8'b00100000;
		color_arr[13597] = 8'b00100000;
		color_arr[13598] = 8'b00100000;
		color_arr[13599] = 8'b00100000;
		color_arr[13600] = 8'b00100000;
		color_arr[13601] = 8'b00100000;
		color_arr[13602] = 8'b00100000;
		color_arr[13603] = 8'b00100000;
		color_arr[13604] = 8'b00100000;
		color_arr[13605] = 8'b00100000;
		color_arr[13606] = 8'b00100000;
		color_arr[13607] = 8'b00100000;
		color_arr[13608] = 8'b00100000;
		color_arr[13609] = 8'b00100000;
		color_arr[13610] = 8'b00100000;
		color_arr[13611] = 8'b00100000;
		color_arr[13612] = 8'b00000000;
		color_arr[13613] = 8'b00000000;
		color_arr[13614] = 8'b00000000;
		color_arr[13615] = 8'b00000000;
		color_arr[13616] = 8'b00000000;
		color_arr[13617] = 8'b00000000;
		color_arr[13618] = 8'b00100000;
		color_arr[13619] = 8'b00100000;
		color_arr[13620] = 8'b00100000;
		color_arr[13621] = 8'b00100000;
		color_arr[13622] = 8'b00100000;
		color_arr[13623] = 8'b00100000;
		color_arr[13624] = 8'b00100000;
		color_arr[13625] = 8'b00100000;
		color_arr[13626] = 8'b00100000;
		color_arr[13627] = 8'b00100000;
		color_arr[13628] = 8'b00100000;
		color_arr[13629] = 8'b00100000;
		color_arr[13630] = 8'b00100000;
		color_arr[13631] = 8'b00100000;
		color_arr[13632] = 8'b00100000;
		color_arr[13633] = 8'b00100000;
		color_arr[13634] = 8'b00100000;
		color_arr[13635] = 8'b00100000;
		color_arr[13636] = 8'b00100000;
		color_arr[13637] = 8'b00100000;
		color_arr[13638] = 8'b00100000;
		color_arr[13639] = 8'b00100000;
		color_arr[13640] = 8'b00100000;
		color_arr[13641] = 8'b00100000;
		color_arr[13642] = 8'b00100000;
		color_arr[13643] = 8'b00100000;
		color_arr[13644] = 8'b00000000;
		color_arr[13645] = 8'b00000000;
		color_arr[13646] = 8'b00000000;
		color_arr[13647] = 8'b00000000;
		color_arr[13648] = 8'b00100000;
		color_arr[13649] = 8'b00100000;
		color_arr[13650] = 8'b00100000;
		color_arr[13651] = 8'b00100000;
		color_arr[13652] = 8'b00100000;
		color_arr[13653] = 8'b00100000;
		color_arr[13654] = 8'b00100000;
		color_arr[13655] = 8'b00100000;
		color_arr[13656] = 8'b00100000;
		color_arr[13657] = 8'b00100000;
		color_arr[13658] = 8'b00100000;
		color_arr[13659] = 8'b00100000;
		color_arr[13660] = 8'b00100000;
		color_arr[13661] = 8'b00000000;
		color_arr[13662] = 8'b00000000;
		color_arr[13663] = 8'b00000000;
		color_arr[13664] = 8'b00000000;
		color_arr[13665] = 8'b00000000;
		color_arr[13666] = 8'b00000000;
		color_arr[13667] = 8'b00100000;
		color_arr[13668] = 8'b00100000;
		color_arr[13669] = 8'b00100000;
		color_arr[13670] = 8'b00100000;
		color_arr[13671] = 8'b00100000;
		color_arr[13672] = 8'b00100000;
		color_arr[13673] = 8'b00100000;
		color_arr[13674] = 8'b00100000;
		color_arr[13675] = 8'b00100000;
		color_arr[13676] = 8'b00100000;
		color_arr[13677] = 8'b00100000;
		color_arr[13678] = 8'b00100000;
		color_arr[13679] = 8'b00100000;
		color_arr[13680] = 8'b00100000;
		color_arr[13681] = 8'b00100000;
		color_arr[13682] = 8'b00100000;
		color_arr[13683] = 8'b00100000;
		color_arr[13684] = 8'b00100000;
		color_arr[13685] = 8'b00100000;
		color_arr[13686] = 8'b00100000;
		color_arr[13687] = 8'b00100000;
		color_arr[13688] = 8'b00000000;
		color_arr[13689] = 8'b00000000;
		color_arr[13690] = 8'b00100000;
		color_arr[13691] = 8'b00100000;
		color_arr[13692] = 8'b00100000;
		color_arr[13693] = 8'b00010010;
		color_arr[13694] = 8'b00010010;
		color_arr[13695] = 8'b00010010;
		color_arr[13696] = 8'b00010010;
		color_arr[13697] = 8'b00010010;
		color_arr[13698] = 8'b00010010;
		color_arr[13699] = 8'b00010010;
		color_arr[13700] = 8'b00010010;
		color_arr[13701] = 8'b00010010;
		color_arr[13702] = 8'b00010010;
		color_arr[13703] = 8'b00010010;
		color_arr[13704] = 8'b00010010;
		color_arr[13705] = 8'b00010010;
		color_arr[13706] = 8'b00010010;
		color_arr[13707] = 8'b00010010;
		color_arr[13708] = 8'b00010010;
		color_arr[13709] = 8'b00010010;
		color_arr[13710] = 8'b00010010;
		color_arr[13711] = 8'b00010010;
		color_arr[13712] = 8'b00010010;
		color_arr[13713] = 8'b00010010;
		color_arr[13714] = 8'b00100000;
		color_arr[13715] = 8'b00100000;
		color_arr[13716] = 8'b00100000;
		color_arr[13717] = 8'b00100000;
		color_arr[13718] = 8'b00100000;
		color_arr[13719] = 8'b00100000;
		color_arr[13720] = 8'b00100000;
		color_arr[13721] = 8'b00100000;
		color_arr[13722] = 8'b00100000;
		color_arr[13723] = 8'b00100000;
		color_arr[13724] = 8'b00100000;
		color_arr[13725] = 8'b00100000;
		color_arr[13726] = 8'b00100000;
		color_arr[13727] = 8'b00100000;
		color_arr[13728] = 8'b00100000;
		color_arr[13729] = 8'b00100000;
		color_arr[13730] = 8'b00100000;
		color_arr[13731] = 8'b00100000;
		color_arr[13732] = 8'b00100000;
		color_arr[13733] = 8'b00100000;
		color_arr[13734] = 8'b00100000;
		color_arr[13735] = 8'b00100000;
		color_arr[13736] = 8'b00100000;
		color_arr[13737] = 8'b00100000;
		color_arr[13738] = 8'b00100000;
		color_arr[13739] = 8'b00000000;
		color_arr[13740] = 8'b00000000;
		color_arr[13741] = 8'b00000000;
		color_arr[13742] = 8'b00000000;
		color_arr[13743] = 8'b00000000;
		color_arr[13744] = 8'b00000000;
		color_arr[13745] = 8'b00100000;
		color_arr[13746] = 8'b00100000;
		color_arr[13747] = 8'b00100000;
		color_arr[13748] = 8'b00100000;
		color_arr[13749] = 8'b00100000;
		color_arr[13750] = 8'b00100000;
		color_arr[13751] = 8'b00100000;
		color_arr[13752] = 8'b00100000;
		color_arr[13753] = 8'b00100000;
		color_arr[13754] = 8'b00100000;
		color_arr[13755] = 8'b00100000;
		color_arr[13756] = 8'b00100000;
		color_arr[13757] = 8'b00100000;
		color_arr[13758] = 8'b00100000;
		color_arr[13759] = 8'b00100000;
		color_arr[13760] = 8'b00100000;
		color_arr[13761] = 8'b00100000;
		color_arr[13762] = 8'b00100000;
		color_arr[13763] = 8'b00100000;
		color_arr[13764] = 8'b00100000;
		color_arr[13765] = 8'b00100000;
		color_arr[13766] = 8'b00100000;
		color_arr[13767] = 8'b00100000;
		color_arr[13768] = 8'b00100000;
		color_arr[13769] = 8'b00100000;
		color_arr[13770] = 8'b00100000;
		color_arr[13771] = 8'b00100000;
		color_arr[13772] = 8'b00100000;
		color_arr[13773] = 8'b00000000;
		color_arr[13774] = 8'b00000000;
		color_arr[13775] = 8'b00000000;
		color_arr[13776] = 8'b00000000;
		color_arr[13777] = 8'b00000000;
		color_arr[13778] = 8'b00000000;
		color_arr[13779] = 8'b00100000;
		color_arr[13780] = 8'b00100000;
		color_arr[13781] = 8'b00100000;
		color_arr[13782] = 8'b00100000;
		color_arr[13783] = 8'b00100000;
		color_arr[13784] = 8'b00100000;
		color_arr[13785] = 8'b00100000;
		color_arr[13786] = 8'b00000000;
		color_arr[13787] = 8'b00000000;
		color_arr[13788] = 8'b00000000;
		color_arr[13789] = 8'b00000000;
		color_arr[13790] = 8'b00000000;
		color_arr[13791] = 8'b00000000;
		color_arr[13792] = 8'b00000000;
		color_arr[13793] = 8'b00100000;
		color_arr[13794] = 8'b00100000;
		color_arr[13795] = 8'b00100000;
		color_arr[13796] = 8'b00100000;
		color_arr[13797] = 8'b00100000;
		color_arr[13798] = 8'b00100000;
		color_arr[13799] = 8'b00100000;
		color_arr[13800] = 8'b00100000;
		color_arr[13801] = 8'b00100000;
		color_arr[13802] = 8'b00100000;
		color_arr[13803] = 8'b00100000;
		color_arr[13804] = 8'b00100000;
		color_arr[13805] = 8'b00100000;
		color_arr[13806] = 8'b00100000;
		color_arr[13807] = 8'b00100000;
		color_arr[13808] = 8'b00100000;
		color_arr[13809] = 8'b00100000;
		color_arr[13810] = 8'b00100000;
		color_arr[13811] = 8'b00100000;
		color_arr[13812] = 8'b00100000;
		color_arr[13813] = 8'b00100000;
		color_arr[13814] = 8'b00100000;
		color_arr[13815] = 8'b00100000;
		color_arr[13816] = 8'b00000000;
		color_arr[13817] = 8'b00000000;
		color_arr[13818] = 8'b00100000;
		color_arr[13819] = 8'b00100000;
		color_arr[13820] = 8'b00100000;
		color_arr[13821] = 8'b00010010;
		color_arr[13822] = 8'b00010010;
		color_arr[13823] = 8'b00010010;
		color_arr[13824] = 8'b00010010;
		color_arr[13825] = 8'b00010010;
		color_arr[13826] = 8'b00010010;
		color_arr[13827] = 8'b00010010;
		color_arr[13828] = 8'b00010010;
		color_arr[13829] = 8'b00010010;
		color_arr[13830] = 8'b00010010;
		color_arr[13831] = 8'b00010010;
		color_arr[13832] = 8'b00010010;
		color_arr[13833] = 8'b00010010;
		color_arr[13834] = 8'b00010010;
		color_arr[13835] = 8'b00010010;
		color_arr[13836] = 8'b00010010;
		color_arr[13837] = 8'b00010010;
		color_arr[13838] = 8'b00010010;
		color_arr[13839] = 8'b00010010;
		color_arr[13840] = 8'b00010010;
		color_arr[13841] = 8'b00010010;
		color_arr[13842] = 8'b00100000;
		color_arr[13843] = 8'b00100000;
		color_arr[13844] = 8'b00100000;
		color_arr[13845] = 8'b00100000;
		color_arr[13846] = 8'b00100000;
		color_arr[13847] = 8'b00100000;
		color_arr[13848] = 8'b00100000;
		color_arr[13849] = 8'b00100000;
		color_arr[13850] = 8'b00100000;
		color_arr[13851] = 8'b00100000;
		color_arr[13852] = 8'b00100000;
		color_arr[13853] = 8'b00100000;
		color_arr[13854] = 8'b00100000;
		color_arr[13855] = 8'b00100000;
		color_arr[13856] = 8'b00100000;
		color_arr[13857] = 8'b00100000;
		color_arr[13858] = 8'b00100000;
		color_arr[13859] = 8'b00100000;
		color_arr[13860] = 8'b00100000;
		color_arr[13861] = 8'b00100000;
		color_arr[13862] = 8'b00100000;
		color_arr[13863] = 8'b00100000;
		color_arr[13864] = 8'b00100000;
		color_arr[13865] = 8'b00100000;
		color_arr[13866] = 8'b00000000;
		color_arr[13867] = 8'b00000000;
		color_arr[13868] = 8'b00000000;
		color_arr[13869] = 8'b00000000;
		color_arr[13870] = 8'b00000000;
		color_arr[13871] = 8'b00000000;
		color_arr[13872] = 8'b00100000;
		color_arr[13873] = 8'b00100000;
		color_arr[13874] = 8'b00100000;
		color_arr[13875] = 8'b00100000;
		color_arr[13876] = 8'b00100000;
		color_arr[13877] = 8'b00100000;
		color_arr[13878] = 8'b00100000;
		color_arr[13879] = 8'b00100000;
		color_arr[13880] = 8'b00100000;
		color_arr[13881] = 8'b00100000;
		color_arr[13882] = 8'b00100000;
		color_arr[13883] = 8'b00100000;
		color_arr[13884] = 8'b00100000;
		color_arr[13885] = 8'b00100000;
		color_arr[13886] = 8'b00100000;
		color_arr[13887] = 8'b00100000;
		color_arr[13888] = 8'b00100000;
		color_arr[13889] = 8'b00100000;
		color_arr[13890] = 8'b00100000;
		color_arr[13891] = 8'b00100000;
		color_arr[13892] = 8'b00100000;
		color_arr[13893] = 8'b00100000;
		color_arr[13894] = 8'b00100000;
		color_arr[13895] = 8'b00100000;
		color_arr[13896] = 8'b00100000;
		color_arr[13897] = 8'b00100000;
		color_arr[13898] = 8'b00100000;
		color_arr[13899] = 8'b00100000;
		color_arr[13900] = 8'b00100000;
		color_arr[13901] = 8'b00100000;
		color_arr[13902] = 8'b00100000;
		color_arr[13903] = 8'b00000000;
		color_arr[13904] = 8'b00000000;
		color_arr[13905] = 8'b00000000;
		color_arr[13906] = 8'b00000000;
		color_arr[13907] = 8'b00000000;
		color_arr[13908] = 8'b00000000;
		color_arr[13909] = 8'b00000000;
		color_arr[13910] = 8'b00000000;
		color_arr[13911] = 8'b00000000;
		color_arr[13912] = 8'b00000000;
		color_arr[13913] = 8'b00000000;
		color_arr[13914] = 8'b00000000;
		color_arr[13915] = 8'b00000000;
		color_arr[13916] = 8'b00000000;
		color_arr[13917] = 8'b00000000;
		color_arr[13918] = 8'b00100000;
		color_arr[13919] = 8'b00100000;
		color_arr[13920] = 8'b00100000;
		color_arr[13921] = 8'b00100000;
		color_arr[13922] = 8'b00100000;
		color_arr[13923] = 8'b00100000;
		color_arr[13924] = 8'b00100000;
		color_arr[13925] = 8'b00100000;
		color_arr[13926] = 8'b00100000;
		color_arr[13927] = 8'b00100000;
		color_arr[13928] = 8'b00100000;
		color_arr[13929] = 8'b00100000;
		color_arr[13930] = 8'b00100000;
		color_arr[13931] = 8'b00100000;
		color_arr[13932] = 8'b00100000;
		color_arr[13933] = 8'b00100000;
		color_arr[13934] = 8'b00100000;
		color_arr[13935] = 8'b00100000;
		color_arr[13936] = 8'b00100000;
		color_arr[13937] = 8'b00100000;
		color_arr[13938] = 8'b00100000;
		color_arr[13939] = 8'b00100000;
		color_arr[13940] = 8'b00100000;
		color_arr[13941] = 8'b00100000;
		color_arr[13942] = 8'b00100000;
		color_arr[13943] = 8'b00100000;
		color_arr[13944] = 8'b00000000;
		color_arr[13945] = 8'b00000000;
		color_arr[13946] = 8'b00100000;
		color_arr[13947] = 8'b00100000;
		color_arr[13948] = 8'b00100000;
		color_arr[13949] = 8'b00010010;
		color_arr[13950] = 8'b00010010;
		color_arr[13951] = 8'b00010010;
		color_arr[13952] = 8'b00010010;
		color_arr[13953] = 8'b00010010;
		color_arr[13954] = 8'b00010010;
		color_arr[13955] = 8'b00010010;
		color_arr[13956] = 8'b00010010;
		color_arr[13957] = 8'b00010010;
		color_arr[13958] = 8'b00010010;
		color_arr[13959] = 8'b00010010;
		color_arr[13960] = 8'b00010010;
		color_arr[13961] = 8'b00010010;
		color_arr[13962] = 8'b00010010;
		color_arr[13963] = 8'b00010010;
		color_arr[13964] = 8'b00010010;
		color_arr[13965] = 8'b00010010;
		color_arr[13966] = 8'b00010010;
		color_arr[13967] = 8'b00010010;
		color_arr[13968] = 8'b00010010;
		color_arr[13969] = 8'b00010010;
		color_arr[13970] = 8'b00100000;
		color_arr[13971] = 8'b00100000;
		color_arr[13972] = 8'b00100000;
		color_arr[13973] = 8'b00100000;
		color_arr[13974] = 8'b00100000;
		color_arr[13975] = 8'b00100000;
		color_arr[13976] = 8'b00100000;
		color_arr[13977] = 8'b00100000;
		color_arr[13978] = 8'b00100000;
		color_arr[13979] = 8'b00100000;
		color_arr[13980] = 8'b00100000;
		color_arr[13981] = 8'b00100000;
		color_arr[13982] = 8'b00100000;
		color_arr[13983] = 8'b00100000;
		color_arr[13984] = 8'b00100000;
		color_arr[13985] = 8'b00100000;
		color_arr[13986] = 8'b00100000;
		color_arr[13987] = 8'b00100000;
		color_arr[13988] = 8'b00100000;
		color_arr[13989] = 8'b00100000;
		color_arr[13990] = 8'b00100000;
		color_arr[13991] = 8'b00100000;
		color_arr[13992] = 8'b00100000;
		color_arr[13993] = 8'b00000000;
		color_arr[13994] = 8'b00000000;
		color_arr[13995] = 8'b00000000;
		color_arr[13996] = 8'b00000000;
		color_arr[13997] = 8'b00000000;
		color_arr[13998] = 8'b00000000;
		color_arr[13999] = 8'b00100000;
		color_arr[14000] = 8'b00100000;
		color_arr[14001] = 8'b00100000;
		color_arr[14002] = 8'b00100000;
		color_arr[14003] = 8'b00100000;
		color_arr[14004] = 8'b00100000;
		color_arr[14005] = 8'b00100000;
		color_arr[14006] = 8'b00100000;
		color_arr[14007] = 8'b00100000;
		color_arr[14008] = 8'b00100000;
		color_arr[14009] = 8'b00100000;
		color_arr[14010] = 8'b00100000;
		color_arr[14011] = 8'b00100000;
		color_arr[14012] = 8'b00100000;
		color_arr[14013] = 8'b00100000;
		color_arr[14014] = 8'b00100000;
		color_arr[14015] = 8'b00100000;
		color_arr[14016] = 8'b00100000;
		color_arr[14017] = 8'b00100000;
		color_arr[14018] = 8'b00100000;
		color_arr[14019] = 8'b00100000;
		color_arr[14020] = 8'b00100000;
		color_arr[14021] = 8'b00100000;
		color_arr[14022] = 8'b00100000;
		color_arr[14023] = 8'b00100000;
		color_arr[14024] = 8'b00100000;
		color_arr[14025] = 8'b00100000;
		color_arr[14026] = 8'b00100000;
		color_arr[14027] = 8'b00100000;
		color_arr[14028] = 8'b00100000;
		color_arr[14029] = 8'b00100000;
		color_arr[14030] = 8'b00100000;
		color_arr[14031] = 8'b00100000;
		color_arr[14032] = 8'b00100000;
		color_arr[14033] = 8'b00100000;
		color_arr[14034] = 8'b00000000;
		color_arr[14035] = 8'b00000000;
		color_arr[14036] = 8'b00000000;
		color_arr[14037] = 8'b00000000;
		color_arr[14038] = 8'b00000000;
		color_arr[14039] = 8'b00000000;
		color_arr[14040] = 8'b00000000;
		color_arr[14041] = 8'b00000000;
		color_arr[14042] = 8'b00000000;
		color_arr[14043] = 8'b00100000;
		color_arr[14044] = 8'b00100000;
		color_arr[14045] = 8'b00100000;
		color_arr[14046] = 8'b00100000;
		color_arr[14047] = 8'b00100000;
		color_arr[14048] = 8'b00100000;
		color_arr[14049] = 8'b00100000;
		color_arr[14050] = 8'b00100000;
		color_arr[14051] = 8'b00100000;
		color_arr[14052] = 8'b00100000;
		color_arr[14053] = 8'b00100000;
		color_arr[14054] = 8'b00100000;
		color_arr[14055] = 8'b00100000;
		color_arr[14056] = 8'b00100000;
		color_arr[14057] = 8'b00100000;
		color_arr[14058] = 8'b00100000;
		color_arr[14059] = 8'b00100000;
		color_arr[14060] = 8'b00100000;
		color_arr[14061] = 8'b00100000;
		color_arr[14062] = 8'b00100000;
		color_arr[14063] = 8'b00100000;
		color_arr[14064] = 8'b00100000;
		color_arr[14065] = 8'b00100000;
		color_arr[14066] = 8'b00100000;
		color_arr[14067] = 8'b00100000;
		color_arr[14068] = 8'b00100000;
		color_arr[14069] = 8'b00100000;
		color_arr[14070] = 8'b00100000;
		color_arr[14071] = 8'b00100000;
		color_arr[14072] = 8'b00000000;
		color_arr[14073] = 8'b00000000;
		color_arr[14074] = 8'b00100000;
		color_arr[14075] = 8'b00100000;
		color_arr[14076] = 8'b00100000;
		color_arr[14077] = 8'b00010010;
		color_arr[14078] = 8'b00010010;
		color_arr[14079] = 8'b00010010;
		color_arr[14080] = 8'b00010010;
		color_arr[14081] = 8'b00010010;
		color_arr[14082] = 8'b00010010;
		color_arr[14083] = 8'b00010010;
		color_arr[14084] = 8'b00010010;
		color_arr[14085] = 8'b00010010;
		color_arr[14086] = 8'b00010010;
		color_arr[14087] = 8'b00010010;
		color_arr[14088] = 8'b00010010;
		color_arr[14089] = 8'b00010010;
		color_arr[14090] = 8'b00010010;
		color_arr[14091] = 8'b00010010;
		color_arr[14092] = 8'b00010010;
		color_arr[14093] = 8'b00010010;
		color_arr[14094] = 8'b00010010;
		color_arr[14095] = 8'b00010010;
		color_arr[14096] = 8'b00010010;
		color_arr[14097] = 8'b00010010;
		color_arr[14098] = 8'b00100000;
		color_arr[14099] = 8'b00100000;
		color_arr[14100] = 8'b00100000;
		color_arr[14101] = 8'b00100000;
		color_arr[14102] = 8'b00100000;
		color_arr[14103] = 8'b00100000;
		color_arr[14104] = 8'b00100000;
		color_arr[14105] = 8'b00100000;
		color_arr[14106] = 8'b00100000;
		color_arr[14107] = 8'b00100000;
		color_arr[14108] = 8'b00100000;
		color_arr[14109] = 8'b00100000;
		color_arr[14110] = 8'b00100000;
		color_arr[14111] = 8'b00100000;
		color_arr[14112] = 8'b00100000;
		color_arr[14113] = 8'b00100000;
		color_arr[14114] = 8'b00100000;
		color_arr[14115] = 8'b00100000;
		color_arr[14116] = 8'b00100000;
		color_arr[14117] = 8'b00100000;
		color_arr[14118] = 8'b00100000;
		color_arr[14119] = 8'b00100000;
		color_arr[14120] = 8'b00000000;
		color_arr[14121] = 8'b00000000;
		color_arr[14122] = 8'b00000000;
		color_arr[14123] = 8'b00000000;
		color_arr[14124] = 8'b00000000;
		color_arr[14125] = 8'b00100000;
		color_arr[14126] = 8'b00100000;
		color_arr[14127] = 8'b00100000;
		color_arr[14128] = 8'b00100000;
		color_arr[14129] = 8'b00100000;
		color_arr[14130] = 8'b00100000;
		color_arr[14131] = 8'b00100000;
		color_arr[14132] = 8'b00100000;
		color_arr[14133] = 8'b00100000;
		color_arr[14134] = 8'b00100000;
		color_arr[14135] = 8'b00100000;
		color_arr[14136] = 8'b00100000;
		color_arr[14137] = 8'b00100000;
		color_arr[14138] = 8'b00100000;
		color_arr[14139] = 8'b00100000;
		color_arr[14140] = 8'b00100000;
		color_arr[14141] = 8'b00100000;
		color_arr[14142] = 8'b00100000;
		color_arr[14143] = 8'b00100000;
		color_arr[14144] = 8'b00100000;
		color_arr[14145] = 8'b00100000;
		color_arr[14146] = 8'b00100000;
		color_arr[14147] = 8'b00100000;
		color_arr[14148] = 8'b00100000;
		color_arr[14149] = 8'b00100000;
		color_arr[14150] = 8'b00100000;
		color_arr[14151] = 8'b00100000;
		color_arr[14152] = 8'b00100000;
		color_arr[14153] = 8'b00100000;
		color_arr[14154] = 8'b00000000;
		color_arr[14155] = 8'b00000000;
		color_arr[14156] = 8'b00000000;
		color_arr[14157] = 8'b00000000;
		color_arr[14158] = 8'b00000000;
		color_arr[14159] = 8'b00000000;
		color_arr[14160] = 8'b00000000;
		color_arr[14161] = 8'b00000000;
		color_arr[14162] = 8'b00000000;
		color_arr[14163] = 8'b00000000;
		color_arr[14164] = 8'b00000000;
		color_arr[14165] = 8'b00000000;
		color_arr[14166] = 8'b00100000;
		color_arr[14167] = 8'b00100000;
		color_arr[14168] = 8'b00100000;
		color_arr[14169] = 8'b00100000;
		color_arr[14170] = 8'b00100000;
		color_arr[14171] = 8'b00100000;
		color_arr[14172] = 8'b00100000;
		color_arr[14173] = 8'b00100000;
		color_arr[14174] = 8'b00100000;
		color_arr[14175] = 8'b00100000;
		color_arr[14176] = 8'b00100000;
		color_arr[14177] = 8'b00100000;
		color_arr[14178] = 8'b00100000;
		color_arr[14179] = 8'b00100000;
		color_arr[14180] = 8'b00100000;
		color_arr[14181] = 8'b00100000;
		color_arr[14182] = 8'b00100000;
		color_arr[14183] = 8'b00100000;
		color_arr[14184] = 8'b00100000;
		color_arr[14185] = 8'b00100000;
		color_arr[14186] = 8'b00100000;
		color_arr[14187] = 8'b00100000;
		color_arr[14188] = 8'b00100000;
		color_arr[14189] = 8'b00100000;
		color_arr[14190] = 8'b00100000;
		color_arr[14191] = 8'b00100000;
		color_arr[14192] = 8'b00100000;
		color_arr[14193] = 8'b00100000;
		color_arr[14194] = 8'b00100000;
		color_arr[14195] = 8'b00100000;
		color_arr[14196] = 8'b00100000;
		color_arr[14197] = 8'b00100000;
		color_arr[14198] = 8'b00100000;
		color_arr[14199] = 8'b00100000;
		color_arr[14200] = 8'b00000000;
		color_arr[14201] = 8'b00000000;
		color_arr[14202] = 8'b00100000;
		color_arr[14203] = 8'b00100000;
		color_arr[14204] = 8'b00100000;
		color_arr[14205] = 8'b00010010;
		color_arr[14206] = 8'b00010010;
		color_arr[14207] = 8'b00010010;
		color_arr[14208] = 8'b00010010;
		color_arr[14209] = 8'b00010010;
		color_arr[14210] = 8'b00010010;
		color_arr[14211] = 8'b00010010;
		color_arr[14212] = 8'b00010010;
		color_arr[14213] = 8'b00010010;
		color_arr[14214] = 8'b00010010;
		color_arr[14215] = 8'b00010010;
		color_arr[14216] = 8'b00010010;
		color_arr[14217] = 8'b00010010;
		color_arr[14218] = 8'b00010010;
		color_arr[14219] = 8'b00010010;
		color_arr[14220] = 8'b00010010;
		color_arr[14221] = 8'b00010010;
		color_arr[14222] = 8'b00010010;
		color_arr[14223] = 8'b00010010;
		color_arr[14224] = 8'b00010010;
		color_arr[14225] = 8'b00010010;
		color_arr[14226] = 8'b00100000;
		color_arr[14227] = 8'b00100000;
		color_arr[14228] = 8'b00100000;
		color_arr[14229] = 8'b00100000;
		color_arr[14230] = 8'b00100000;
		color_arr[14231] = 8'b00100000;
		color_arr[14232] = 8'b00100000;
		color_arr[14233] = 8'b00100000;
		color_arr[14234] = 8'b00100000;
		color_arr[14235] = 8'b00100000;
		color_arr[14236] = 8'b00100000;
		color_arr[14237] = 8'b00100000;
		color_arr[14238] = 8'b00100000;
		color_arr[14239] = 8'b00100000;
		color_arr[14240] = 8'b00100000;
		color_arr[14241] = 8'b00100000;
		color_arr[14242] = 8'b00100000;
		color_arr[14243] = 8'b00100000;
		color_arr[14244] = 8'b00100000;
		color_arr[14245] = 8'b00100000;
		color_arr[14246] = 8'b00100000;
		color_arr[14247] = 8'b00000000;
		color_arr[14248] = 8'b00000000;
		color_arr[14249] = 8'b00000000;
		color_arr[14250] = 8'b00000000;
		color_arr[14251] = 8'b00000000;
		color_arr[14252] = 8'b00100000;
		color_arr[14253] = 8'b00100000;
		color_arr[14254] = 8'b00100000;
		color_arr[14255] = 8'b00100000;
		color_arr[14256] = 8'b00100000;
		color_arr[14257] = 8'b00100000;
		color_arr[14258] = 8'b00100000;
		color_arr[14259] = 8'b00100000;
		color_arr[14260] = 8'b00100000;
		color_arr[14261] = 8'b00100000;
		color_arr[14262] = 8'b00100000;
		color_arr[14263] = 8'b00100000;
		color_arr[14264] = 8'b00100000;
		color_arr[14265] = 8'b00100000;
		color_arr[14266] = 8'b00100000;
		color_arr[14267] = 8'b00100000;
		color_arr[14268] = 8'b00100000;
		color_arr[14269] = 8'b00100000;
		color_arr[14270] = 8'b00100000;
		color_arr[14271] = 8'b00100000;
		color_arr[14272] = 8'b00100000;
		color_arr[14273] = 8'b00100000;
		color_arr[14274] = 8'b00100000;
		color_arr[14275] = 8'b00100000;
		color_arr[14276] = 8'b00000000;
		color_arr[14277] = 8'b00000000;
		color_arr[14278] = 8'b00000000;
		color_arr[14279] = 8'b00000000;
		color_arr[14280] = 8'b00000000;
		color_arr[14281] = 8'b00000000;
		color_arr[14282] = 8'b00000000;
		color_arr[14283] = 8'b00000000;
		color_arr[14284] = 8'b00000000;
		color_arr[14285] = 8'b00000000;
		color_arr[14286] = 8'b00000000;
		color_arr[14287] = 8'b00000000;
		color_arr[14288] = 8'b00000000;
		color_arr[14289] = 8'b00000000;
		color_arr[14290] = 8'b00000000;
		color_arr[14291] = 8'b00000000;
		color_arr[14292] = 8'b00000000;
		color_arr[14293] = 8'b00000000;
		color_arr[14294] = 8'b00000000;
		color_arr[14295] = 8'b00000000;
		color_arr[14296] = 8'b00000000;
		color_arr[14297] = 8'b00000000;
		color_arr[14298] = 8'b00100000;
		color_arr[14299] = 8'b00100000;
		color_arr[14300] = 8'b00100000;
		color_arr[14301] = 8'b00100000;
		color_arr[14302] = 8'b00100000;
		color_arr[14303] = 8'b00100000;
		color_arr[14304] = 8'b00100000;
		color_arr[14305] = 8'b00100000;
		color_arr[14306] = 8'b00100000;
		color_arr[14307] = 8'b00100000;
		color_arr[14308] = 8'b00100000;
		color_arr[14309] = 8'b00100000;
		color_arr[14310] = 8'b00100000;
		color_arr[14311] = 8'b00100000;
		color_arr[14312] = 8'b00100000;
		color_arr[14313] = 8'b00100000;
		color_arr[14314] = 8'b00100000;
		color_arr[14315] = 8'b00100000;
		color_arr[14316] = 8'b00100000;
		color_arr[14317] = 8'b00100000;
		color_arr[14318] = 8'b00100000;
		color_arr[14319] = 8'b00100000;
		color_arr[14320] = 8'b00100000;
		color_arr[14321] = 8'b00100000;
		color_arr[14322] = 8'b00100000;
		color_arr[14323] = 8'b00100000;
		color_arr[14324] = 8'b00100000;
		color_arr[14325] = 8'b00100000;
		color_arr[14326] = 8'b00100000;
		color_arr[14327] = 8'b00100000;
		color_arr[14328] = 8'b00000000;
		color_arr[14329] = 8'b00000000;
		color_arr[14330] = 8'b00000000;
		color_arr[14331] = 8'b00100000;
		color_arr[14332] = 8'b00100000;
		color_arr[14333] = 8'b00010010;
		color_arr[14334] = 8'b00010010;
		color_arr[14335] = 8'b00010010;
		color_arr[14336] = 8'b00000000;
		color_arr[14337] = 8'b00010010;
		color_arr[14338] = 8'b00010010;
		color_arr[14339] = 8'b00010010;
		color_arr[14340] = 8'b00010010;
		color_arr[14341] = 8'b00010010;
		color_arr[14342] = 8'b00010010;
		color_arr[14343] = 8'b00010010;
		color_arr[14344] = 8'b00010010;
		color_arr[14345] = 8'b00010010;
		color_arr[14346] = 8'b00010010;
		color_arr[14347] = 8'b00010010;
		color_arr[14348] = 8'b00010010;
		color_arr[14349] = 8'b00010010;
		color_arr[14350] = 8'b00010010;
		color_arr[14351] = 8'b00010010;
		color_arr[14352] = 8'b00010010;
		color_arr[14353] = 8'b00010010;
		color_arr[14354] = 8'b00100000;
		color_arr[14355] = 8'b00100000;
		color_arr[14356] = 8'b00100000;
		color_arr[14357] = 8'b00100000;
		color_arr[14358] = 8'b00100000;
		color_arr[14359] = 8'b00100000;
		color_arr[14360] = 8'b00100000;
		color_arr[14361] = 8'b00100000;
		color_arr[14362] = 8'b00100000;
		color_arr[14363] = 8'b00100000;
		color_arr[14364] = 8'b00100000;
		color_arr[14365] = 8'b00100000;
		color_arr[14366] = 8'b00100000;
		color_arr[14367] = 8'b00100000;
		color_arr[14368] = 8'b00100000;
		color_arr[14369] = 8'b00100000;
		color_arr[14370] = 8'b00100000;
		color_arr[14371] = 8'b00100000;
		color_arr[14372] = 8'b00100000;
		color_arr[14373] = 8'b00100000;
		color_arr[14374] = 8'b00000000;
		color_arr[14375] = 8'b00000000;
		color_arr[14376] = 8'b00000000;
		color_arr[14377] = 8'b00000000;
		color_arr[14378] = 8'b00000000;
		color_arr[14379] = 8'b00100000;
		color_arr[14380] = 8'b00100000;
		color_arr[14381] = 8'b00100000;
		color_arr[14382] = 8'b00100000;
		color_arr[14383] = 8'b00100000;
		color_arr[14384] = 8'b00100000;
		color_arr[14385] = 8'b00100000;
		color_arr[14386] = 8'b00100000;
		color_arr[14387] = 8'b00100000;
		color_arr[14388] = 8'b00100000;
		color_arr[14389] = 8'b00100000;
		color_arr[14390] = 8'b00100000;
		color_arr[14391] = 8'b00100000;
		color_arr[14392] = 8'b00100000;
		color_arr[14393] = 8'b00100000;
		color_arr[14394] = 8'b00100000;
		color_arr[14395] = 8'b00100000;
		color_arr[14396] = 8'b00100000;
		color_arr[14397] = 8'b00100000;
		color_arr[14398] = 8'b00100000;
		color_arr[14399] = 8'b00100000;
		color_arr[14400] = 8'b00000000;
		color_arr[14401] = 8'b00000000;
		color_arr[14402] = 8'b00000000;
		color_arr[14403] = 8'b00000000;
		color_arr[14404] = 8'b00000000;
		color_arr[14405] = 8'b00000000;
		color_arr[14406] = 8'b00000000;
		color_arr[14407] = 8'b00000000;
		color_arr[14408] = 8'b00000000;
		color_arr[14409] = 8'b00000000;
		color_arr[14410] = 8'b00000000;
		color_arr[14411] = 8'b00100000;
		color_arr[14412] = 8'b00100000;
		color_arr[14413] = 8'b00100000;
		color_arr[14414] = 8'b00100000;
		color_arr[14415] = 8'b00100000;
		color_arr[14416] = 8'b00100000;
		color_arr[14417] = 8'b00100000;
		color_arr[14418] = 8'b00100000;
		color_arr[14419] = 8'b00100000;
		color_arr[14420] = 8'b00100000;
		color_arr[14421] = 8'b00000000;
		color_arr[14422] = 8'b00000000;
		color_arr[14423] = 8'b00000000;
		color_arr[14424] = 8'b00000000;
		color_arr[14425] = 8'b00000000;
		color_arr[14426] = 8'b00000000;
		color_arr[14427] = 8'b00000000;
		color_arr[14428] = 8'b00000000;
		color_arr[14429] = 8'b00000000;
		color_arr[14430] = 8'b00100000;
		color_arr[14431] = 8'b00100000;
		color_arr[14432] = 8'b00100000;
		color_arr[14433] = 8'b00100000;
		color_arr[14434] = 8'b00100000;
		color_arr[14435] = 8'b00100000;
		color_arr[14436] = 8'b00100000;
		color_arr[14437] = 8'b00100000;
		color_arr[14438] = 8'b00100000;
		color_arr[14439] = 8'b00100000;
		color_arr[14440] = 8'b00100000;
		color_arr[14441] = 8'b00100000;
		color_arr[14442] = 8'b00100000;
		color_arr[14443] = 8'b00100000;
		color_arr[14444] = 8'b00100000;
		color_arr[14445] = 8'b00100000;
		color_arr[14446] = 8'b00100000;
		color_arr[14447] = 8'b00100000;
		color_arr[14448] = 8'b00100000;
		color_arr[14449] = 8'b00100000;
		color_arr[14450] = 8'b00100000;
		color_arr[14451] = 8'b00100000;
		color_arr[14452] = 8'b00100000;
		color_arr[14453] = 8'b00100000;
		color_arr[14454] = 8'b00100000;
		color_arr[14455] = 8'b00100000;
		color_arr[14456] = 8'b00100000;
		color_arr[14457] = 8'b00000000;
		color_arr[14458] = 8'b00000000;
		color_arr[14459] = 8'b00100000;
		color_arr[14460] = 8'b00100000;
		color_arr[14461] = 8'b00010010;
		color_arr[14462] = 8'b00010010;
		color_arr[14463] = 8'b00010010;
		color_arr[14464] = 8'b00000000;
		color_arr[14465] = 8'b00010010;
		color_arr[14466] = 8'b00010010;
		color_arr[14467] = 8'b00010010;
		color_arr[14468] = 8'b00010010;
		color_arr[14469] = 8'b00010010;
		color_arr[14470] = 8'b00010010;
		color_arr[14471] = 8'b00010010;
		color_arr[14472] = 8'b00010010;
		color_arr[14473] = 8'b00010010;
		color_arr[14474] = 8'b00010010;
		color_arr[14475] = 8'b00010010;
		color_arr[14476] = 8'b00010010;
		color_arr[14477] = 8'b00010010;
		color_arr[14478] = 8'b00010010;
		color_arr[14479] = 8'b00010010;
		color_arr[14480] = 8'b00010010;
		color_arr[14481] = 8'b00010010;
		color_arr[14482] = 8'b00100000;
		color_arr[14483] = 8'b00100000;
		color_arr[14484] = 8'b00100000;
		color_arr[14485] = 8'b00100000;
		color_arr[14486] = 8'b00100000;
		color_arr[14487] = 8'b00100000;
		color_arr[14488] = 8'b00100000;
		color_arr[14489] = 8'b00100000;
		color_arr[14490] = 8'b00100000;
		color_arr[14491] = 8'b00100000;
		color_arr[14492] = 8'b00100000;
		color_arr[14493] = 8'b00100000;
		color_arr[14494] = 8'b00100000;
		color_arr[14495] = 8'b00100000;
		color_arr[14496] = 8'b00100000;
		color_arr[14497] = 8'b00100000;
		color_arr[14498] = 8'b00100000;
		color_arr[14499] = 8'b00100000;
		color_arr[14500] = 8'b00100000;
		color_arr[14501] = 8'b00000000;
		color_arr[14502] = 8'b00000000;
		color_arr[14503] = 8'b00000000;
		color_arr[14504] = 8'b00000000;
		color_arr[14505] = 8'b00000000;
		color_arr[14506] = 8'b00100000;
		color_arr[14507] = 8'b00100000;
		color_arr[14508] = 8'b00100000;
		color_arr[14509] = 8'b00100000;
		color_arr[14510] = 8'b00100000;
		color_arr[14511] = 8'b00100000;
		color_arr[14512] = 8'b00100000;
		color_arr[14513] = 8'b00100000;
		color_arr[14514] = 8'b00100000;
		color_arr[14515] = 8'b00100000;
		color_arr[14516] = 8'b00100000;
		color_arr[14517] = 8'b00100000;
		color_arr[14518] = 8'b00100000;
		color_arr[14519] = 8'b00100000;
		color_arr[14520] = 8'b00100000;
		color_arr[14521] = 8'b00100000;
		color_arr[14522] = 8'b00100000;
		color_arr[14523] = 8'b00100000;
		color_arr[14524] = 8'b00100000;
		color_arr[14525] = 8'b00000000;
		color_arr[14526] = 8'b00000000;
		color_arr[14527] = 8'b00000000;
		color_arr[14528] = 8'b00000000;
		color_arr[14529] = 8'b00000000;
		color_arr[14530] = 8'b00000000;
		color_arr[14531] = 8'b00000000;
		color_arr[14532] = 8'b00000000;
		color_arr[14533] = 8'b00100000;
		color_arr[14534] = 8'b00100000;
		color_arr[14535] = 8'b00100000;
		color_arr[14536] = 8'b00100000;
		color_arr[14537] = 8'b00100000;
		color_arr[14538] = 8'b00100000;
		color_arr[14539] = 8'b00100000;
		color_arr[14540] = 8'b00100000;
		color_arr[14541] = 8'b00100000;
		color_arr[14542] = 8'b00100000;
		color_arr[14543] = 8'b00100000;
		color_arr[14544] = 8'b00100000;
		color_arr[14545] = 8'b00100000;
		color_arr[14546] = 8'b00100000;
		color_arr[14547] = 8'b00100000;
		color_arr[14548] = 8'b00100000;
		color_arr[14549] = 8'b00100000;
		color_arr[14550] = 8'b00100000;
		color_arr[14551] = 8'b00100000;
		color_arr[14552] = 8'b00100000;
		color_arr[14553] = 8'b00000000;
		color_arr[14554] = 8'b00000000;
		color_arr[14555] = 8'b00000000;
		color_arr[14556] = 8'b00000000;
		color_arr[14557] = 8'b00000000;
		color_arr[14558] = 8'b00000000;
		color_arr[14559] = 8'b00000000;
		color_arr[14560] = 8'b00000000;
		color_arr[14561] = 8'b00000000;
		color_arr[14562] = 8'b00100000;
		color_arr[14563] = 8'b00100000;
		color_arr[14564] = 8'b00100000;
		color_arr[14565] = 8'b00100000;
		color_arr[14566] = 8'b00100000;
		color_arr[14567] = 8'b00100000;
		color_arr[14568] = 8'b00100000;
		color_arr[14569] = 8'b00100000;
		color_arr[14570] = 8'b00100000;
		color_arr[14571] = 8'b00100000;
		color_arr[14572] = 8'b00100000;
		color_arr[14573] = 8'b00100000;
		color_arr[14574] = 8'b00100000;
		color_arr[14575] = 8'b00100000;
		color_arr[14576] = 8'b00100000;
		color_arr[14577] = 8'b00100000;
		color_arr[14578] = 8'b00100000;
		color_arr[14579] = 8'b00100000;
		color_arr[14580] = 8'b00100000;
		color_arr[14581] = 8'b00100000;
		color_arr[14582] = 8'b00100000;
		color_arr[14583] = 8'b00100000;
		color_arr[14584] = 8'b00100000;
		color_arr[14585] = 8'b00000000;
		color_arr[14586] = 8'b00000000;
		color_arr[14587] = 8'b00100000;
		color_arr[14588] = 8'b00100000;
		color_arr[14589] = 8'b00010010;
		color_arr[14590] = 8'b00010010;
		color_arr[14591] = 8'b00010010;
		color_arr[14592] = 8'b00000000;
		color_arr[14593] = 8'b00000000;
		color_arr[14594] = 8'b00010010;
		color_arr[14595] = 8'b00010010;
		color_arr[14596] = 8'b00010010;
		color_arr[14597] = 8'b00010010;
		color_arr[14598] = 8'b00010010;
		color_arr[14599] = 8'b00010010;
		color_arr[14600] = 8'b00010010;
		color_arr[14601] = 8'b00010010;
		color_arr[14602] = 8'b00010010;
		color_arr[14603] = 8'b00010010;
		color_arr[14604] = 8'b00010010;
		color_arr[14605] = 8'b00010010;
		color_arr[14606] = 8'b00010010;
		color_arr[14607] = 8'b00010010;
		color_arr[14608] = 8'b00010010;
		color_arr[14609] = 8'b00010010;
		color_arr[14610] = 8'b00100000;
		color_arr[14611] = 8'b00100000;
		color_arr[14612] = 8'b00100000;
		color_arr[14613] = 8'b00100000;
		color_arr[14614] = 8'b00100000;
		color_arr[14615] = 8'b00100000;
		color_arr[14616] = 8'b00100000;
		color_arr[14617] = 8'b00100000;
		color_arr[14618] = 8'b00100000;
		color_arr[14619] = 8'b00100000;
		color_arr[14620] = 8'b00100000;
		color_arr[14621] = 8'b00100000;
		color_arr[14622] = 8'b00100000;
		color_arr[14623] = 8'b00100000;
		color_arr[14624] = 8'b00100000;
		color_arr[14625] = 8'b00100000;
		color_arr[14626] = 8'b00100000;
		color_arr[14627] = 8'b00100000;
		color_arr[14628] = 8'b00000000;
		color_arr[14629] = 8'b00000000;
		color_arr[14630] = 8'b00000000;
		color_arr[14631] = 8'b00000000;
		color_arr[14632] = 8'b00000000;
		color_arr[14633] = 8'b00100000;
		color_arr[14634] = 8'b00100000;
		color_arr[14635] = 8'b00100000;
		color_arr[14636] = 8'b00100000;
		color_arr[14637] = 8'b00100000;
		color_arr[14638] = 8'b00100000;
		color_arr[14639] = 8'b00100000;
		color_arr[14640] = 8'b00100000;
		color_arr[14641] = 8'b00100000;
		color_arr[14642] = 8'b00100000;
		color_arr[14643] = 8'b00100000;
		color_arr[14644] = 8'b00100000;
		color_arr[14645] = 8'b00100000;
		color_arr[14646] = 8'b00100000;
		color_arr[14647] = 8'b00100000;
		color_arr[14648] = 8'b00100000;
		color_arr[14649] = 8'b00100000;
		color_arr[14650] = 8'b00000000;
		color_arr[14651] = 8'b00000000;
		color_arr[14652] = 8'b00000000;
		color_arr[14653] = 8'b00000000;
		color_arr[14654] = 8'b00000000;
		color_arr[14655] = 8'b00000000;
		color_arr[14656] = 8'b00000000;
		color_arr[14657] = 8'b00100000;
		color_arr[14658] = 8'b00100000;
		color_arr[14659] = 8'b00100000;
		color_arr[14660] = 8'b00100000;
		color_arr[14661] = 8'b00100000;
		color_arr[14662] = 8'b00100000;
		color_arr[14663] = 8'b00100000;
		color_arr[14664] = 8'b00100000;
		color_arr[14665] = 8'b00100000;
		color_arr[14666] = 8'b00100000;
		color_arr[14667] = 8'b00100000;
		color_arr[14668] = 8'b00100000;
		color_arr[14669] = 8'b00100000;
		color_arr[14670] = 8'b00100000;
		color_arr[14671] = 8'b00100000;
		color_arr[14672] = 8'b00100000;
		color_arr[14673] = 8'b00100000;
		color_arr[14674] = 8'b00100000;
		color_arr[14675] = 8'b00100000;
		color_arr[14676] = 8'b00100000;
		color_arr[14677] = 8'b00100000;
		color_arr[14678] = 8'b00100000;
		color_arr[14679] = 8'b00100000;
		color_arr[14680] = 8'b00100000;
		color_arr[14681] = 8'b00100000;
		color_arr[14682] = 8'b00100000;
		color_arr[14683] = 8'b00100000;
		color_arr[14684] = 8'b00100000;
		color_arr[14685] = 8'b00000000;
		color_arr[14686] = 8'b00000000;
		color_arr[14687] = 8'b00000000;
		color_arr[14688] = 8'b00000000;
		color_arr[14689] = 8'b00000000;
		color_arr[14690] = 8'b00000000;
		color_arr[14691] = 8'b00000000;
		color_arr[14692] = 8'b00000000;
		color_arr[14693] = 8'b00000000;
		color_arr[14694] = 8'b00100000;
		color_arr[14695] = 8'b00100000;
		color_arr[14696] = 8'b00100000;
		color_arr[14697] = 8'b00100000;
		color_arr[14698] = 8'b00100000;
		color_arr[14699] = 8'b00100000;
		color_arr[14700] = 8'b00100000;
		color_arr[14701] = 8'b00100000;
		color_arr[14702] = 8'b00100000;
		color_arr[14703] = 8'b00100000;
		color_arr[14704] = 8'b00100000;
		color_arr[14705] = 8'b00100000;
		color_arr[14706] = 8'b00100000;
		color_arr[14707] = 8'b00100000;
		color_arr[14708] = 8'b00100000;
		color_arr[14709] = 8'b00100000;
		color_arr[14710] = 8'b00100000;
		color_arr[14711] = 8'b00100000;
		color_arr[14712] = 8'b00100000;
		color_arr[14713] = 8'b00000000;
		color_arr[14714] = 8'b00000000;
		color_arr[14715] = 8'b00100000;
		color_arr[14716] = 8'b00100000;
		color_arr[14717] = 8'b00010010;
		color_arr[14718] = 8'b00010010;
		color_arr[14719] = 8'b00010010;
		color_arr[14720] = 8'b00000000;
		color_arr[14721] = 8'b00000000;
		color_arr[14722] = 8'b00000000;
		color_arr[14723] = 8'b00000000;
		color_arr[14724] = 8'b00010010;
		color_arr[14725] = 8'b00010010;
		color_arr[14726] = 8'b00010010;
		color_arr[14727] = 8'b00010010;
		color_arr[14728] = 8'b00010010;
		color_arr[14729] = 8'b00010010;
		color_arr[14730] = 8'b00010010;
		color_arr[14731] = 8'b00010010;
		color_arr[14732] = 8'b00010010;
		color_arr[14733] = 8'b00010010;
		color_arr[14734] = 8'b00010010;
		color_arr[14735] = 8'b00010010;
		color_arr[14736] = 8'b00010010;
		color_arr[14737] = 8'b00010010;
		color_arr[14738] = 8'b00100000;
		color_arr[14739] = 8'b00100000;
		color_arr[14740] = 8'b00100000;
		color_arr[14741] = 8'b00100000;
		color_arr[14742] = 8'b00100000;
		color_arr[14743] = 8'b00100000;
		color_arr[14744] = 8'b00100000;
		color_arr[14745] = 8'b00100000;
		color_arr[14746] = 8'b00100000;
		color_arr[14747] = 8'b00100000;
		color_arr[14748] = 8'b00100000;
		color_arr[14749] = 8'b00100000;
		color_arr[14750] = 8'b00100000;
		color_arr[14751] = 8'b00100000;
		color_arr[14752] = 8'b00100000;
		color_arr[14753] = 8'b00100000;
		color_arr[14754] = 8'b00100000;
		color_arr[14755] = 8'b00000000;
		color_arr[14756] = 8'b00000000;
		color_arr[14757] = 8'b00000000;
		color_arr[14758] = 8'b00000000;
		color_arr[14759] = 8'b00100000;
		color_arr[14760] = 8'b00100000;
		color_arr[14761] = 8'b00100000;
		color_arr[14762] = 8'b00100000;
		color_arr[14763] = 8'b00100000;
		color_arr[14764] = 8'b00100000;
		color_arr[14765] = 8'b00100000;
		color_arr[14766] = 8'b00100000;
		color_arr[14767] = 8'b00100000;
		color_arr[14768] = 8'b00100000;
		color_arr[14769] = 8'b00100000;
		color_arr[14770] = 8'b00100000;
		color_arr[14771] = 8'b00100000;
		color_arr[14772] = 8'b00100000;
		color_arr[14773] = 8'b00100000;
		color_arr[14774] = 8'b00100000;
		color_arr[14775] = 8'b00000000;
		color_arr[14776] = 8'b00000000;
		color_arr[14777] = 8'b00000000;
		color_arr[14778] = 8'b00000000;
		color_arr[14779] = 8'b00000000;
		color_arr[14780] = 8'b00000000;
		color_arr[14781] = 8'b00000000;
		color_arr[14782] = 8'b00100000;
		color_arr[14783] = 8'b00100000;
		color_arr[14784] = 8'b00100000;
		color_arr[14785] = 8'b00100000;
		color_arr[14786] = 8'b00100000;
		color_arr[14787] = 8'b00100000;
		color_arr[14788] = 8'b00100000;
		color_arr[14789] = 8'b00100000;
		color_arr[14790] = 8'b00100000;
		color_arr[14791] = 8'b00100000;
		color_arr[14792] = 8'b00100000;
		color_arr[14793] = 8'b00100000;
		color_arr[14794] = 8'b00100000;
		color_arr[14795] = 8'b00100000;
		color_arr[14796] = 8'b00100000;
		color_arr[14797] = 8'b00100000;
		color_arr[14798] = 8'b00100000;
		color_arr[14799] = 8'b00100000;
		color_arr[14800] = 8'b00100000;
		color_arr[14801] = 8'b00100000;
		color_arr[14802] = 8'b00100000;
		color_arr[14803] = 8'b00100000;
		color_arr[14804] = 8'b00100000;
		color_arr[14805] = 8'b00100000;
		color_arr[14806] = 8'b00100000;
		color_arr[14807] = 8'b00100000;
		color_arr[14808] = 8'b00100000;
		color_arr[14809] = 8'b00100000;
		color_arr[14810] = 8'b00100000;
		color_arr[14811] = 8'b00100000;
		color_arr[14812] = 8'b00100000;
		color_arr[14813] = 8'b00100000;
		color_arr[14814] = 8'b00100000;
		color_arr[14815] = 8'b00100000;
		color_arr[14816] = 8'b00100000;
		color_arr[14817] = 8'b00000000;
		color_arr[14818] = 8'b00000000;
		color_arr[14819] = 8'b00000000;
		color_arr[14820] = 8'b00000000;
		color_arr[14821] = 8'b00000000;
		color_arr[14822] = 8'b00000000;
		color_arr[14823] = 8'b00000000;
		color_arr[14824] = 8'b00100000;
		color_arr[14825] = 8'b00100000;
		color_arr[14826] = 8'b00100000;
		color_arr[14827] = 8'b00100000;
		color_arr[14828] = 8'b00100000;
		color_arr[14829] = 8'b00100000;
		color_arr[14830] = 8'b00100000;
		color_arr[14831] = 8'b00100000;
		color_arr[14832] = 8'b00100000;
		color_arr[14833] = 8'b00100000;
		color_arr[14834] = 8'b00100000;
		color_arr[14835] = 8'b00100000;
		color_arr[14836] = 8'b00100000;
		color_arr[14837] = 8'b00100000;
		color_arr[14838] = 8'b00100000;
		color_arr[14839] = 8'b00100000;
		color_arr[14840] = 8'b00100000;
		color_arr[14841] = 8'b00000000;
		color_arr[14842] = 8'b00000000;
		color_arr[14843] = 8'b00100000;
		color_arr[14844] = 8'b00100000;
		color_arr[14845] = 8'b00010010;
		color_arr[14846] = 8'b00010010;
		color_arr[14847] = 8'b00010010;
		color_arr[14848] = 8'b00010010;
		color_arr[14849] = 8'b00000000;
		color_arr[14850] = 8'b00000000;
		color_arr[14851] = 8'b00000000;
		color_arr[14852] = 8'b00000000;
		color_arr[14853] = 8'b00010010;
		color_arr[14854] = 8'b00010010;
		color_arr[14855] = 8'b00010010;
		color_arr[14856] = 8'b00010010;
		color_arr[14857] = 8'b00010010;
		color_arr[14858] = 8'b00010010;
		color_arr[14859] = 8'b00010010;
		color_arr[14860] = 8'b00010010;
		color_arr[14861] = 8'b00010010;
		color_arr[14862] = 8'b00010010;
		color_arr[14863] = 8'b00010010;
		color_arr[14864] = 8'b00010010;
		color_arr[14865] = 8'b00010010;
		color_arr[14866] = 8'b00100000;
		color_arr[14867] = 8'b00100000;
		color_arr[14868] = 8'b00100000;
		color_arr[14869] = 8'b00100000;
		color_arr[14870] = 8'b00100000;
		color_arr[14871] = 8'b00100000;
		color_arr[14872] = 8'b00100000;
		color_arr[14873] = 8'b00100000;
		color_arr[14874] = 8'b00100000;
		color_arr[14875] = 8'b00100000;
		color_arr[14876] = 8'b00100000;
		color_arr[14877] = 8'b00100000;
		color_arr[14878] = 8'b00100000;
		color_arr[14879] = 8'b00100000;
		color_arr[14880] = 8'b00100000;
		color_arr[14881] = 8'b00100000;
		color_arr[14882] = 8'b00000000;
		color_arr[14883] = 8'b00000000;
		color_arr[14884] = 8'b00000000;
		color_arr[14885] = 8'b00000000;
		color_arr[14886] = 8'b00100000;
		color_arr[14887] = 8'b00100000;
		color_arr[14888] = 8'b00100000;
		color_arr[14889] = 8'b00100000;
		color_arr[14890] = 8'b00100000;
		color_arr[14891] = 8'b00100000;
		color_arr[14892] = 8'b00100000;
		color_arr[14893] = 8'b00100000;
		color_arr[14894] = 8'b00100000;
		color_arr[14895] = 8'b00100000;
		color_arr[14896] = 8'b00100000;
		color_arr[14897] = 8'b00100000;
		color_arr[14898] = 8'b00100000;
		color_arr[14899] = 8'b00100000;
		color_arr[14900] = 8'b00100000;
		color_arr[14901] = 8'b00000000;
		color_arr[14902] = 8'b00000000;
		color_arr[14903] = 8'b00000000;
		color_arr[14904] = 8'b00000000;
		color_arr[14905] = 8'b00000000;
		color_arr[14906] = 8'b00000000;
		color_arr[14907] = 8'b00100000;
		color_arr[14908] = 8'b00100000;
		color_arr[14909] = 8'b00100000;
		color_arr[14910] = 8'b00100000;
		color_arr[14911] = 8'b00100000;
		color_arr[14912] = 8'b00100000;
		color_arr[14913] = 8'b00100000;
		color_arr[14914] = 8'b00100000;
		color_arr[14915] = 8'b00100000;
		color_arr[14916] = 8'b00100000;
		color_arr[14917] = 8'b00100000;
		color_arr[14918] = 8'b00100000;
		color_arr[14919] = 8'b00100000;
		color_arr[14920] = 8'b00100000;
		color_arr[14921] = 8'b00100000;
		color_arr[14922] = 8'b00100000;
		color_arr[14923] = 8'b00100000;
		color_arr[14924] = 8'b00100000;
		color_arr[14925] = 8'b00100000;
		color_arr[14926] = 8'b00100000;
		color_arr[14927] = 8'b00100000;
		color_arr[14928] = 8'b00100000;
		color_arr[14929] = 8'b00100000;
		color_arr[14930] = 8'b00100000;
		color_arr[14931] = 8'b00100000;
		color_arr[14932] = 8'b00100000;
		color_arr[14933] = 8'b00100000;
		color_arr[14934] = 8'b00100000;
		color_arr[14935] = 8'b00100000;
		color_arr[14936] = 8'b00100000;
		color_arr[14937] = 8'b00100000;
		color_arr[14938] = 8'b00100000;
		color_arr[14939] = 8'b00100000;
		color_arr[14940] = 8'b00100000;
		color_arr[14941] = 8'b00100000;
		color_arr[14942] = 8'b00100000;
		color_arr[14943] = 8'b00100000;
		color_arr[14944] = 8'b00100000;
		color_arr[14945] = 8'b00100000;
		color_arr[14946] = 8'b00100000;
		color_arr[14947] = 8'b00100000;
		color_arr[14948] = 8'b00100000;
		color_arr[14949] = 8'b00000000;
		color_arr[14950] = 8'b00000000;
		color_arr[14951] = 8'b00000000;
		color_arr[14952] = 8'b00000000;
		color_arr[14953] = 8'b00000000;
		color_arr[14954] = 8'b00000000;
		color_arr[14955] = 8'b00100000;
		color_arr[14956] = 8'b00100000;
		color_arr[14957] = 8'b00100000;
		color_arr[14958] = 8'b00100000;
		color_arr[14959] = 8'b00100000;
		color_arr[14960] = 8'b00100000;
		color_arr[14961] = 8'b00100000;
		color_arr[14962] = 8'b00100000;
		color_arr[14963] = 8'b00100000;
		color_arr[14964] = 8'b00100000;
		color_arr[14965] = 8'b00100000;
		color_arr[14966] = 8'b00100000;
		color_arr[14967] = 8'b00100000;
		color_arr[14968] = 8'b00100000;
		color_arr[14969] = 8'b00000000;
		color_arr[14970] = 8'b00000000;
		color_arr[14971] = 8'b00100000;
		color_arr[14972] = 8'b00100000;
		color_arr[14973] = 8'b00010010;
		color_arr[14974] = 8'b00010010;
		color_arr[14975] = 8'b00010010;
		color_arr[14976] = 8'b00010010;
		color_arr[14977] = 8'b00010010;
		color_arr[14978] = 8'b00010010;
		color_arr[14979] = 8'b00000000;
		color_arr[14980] = 8'b00000000;
		color_arr[14981] = 8'b00000000;
		color_arr[14982] = 8'b00000000;
		color_arr[14983] = 8'b00010010;
		color_arr[14984] = 8'b00010010;
		color_arr[14985] = 8'b00010010;
		color_arr[14986] = 8'b00010010;
		color_arr[14987] = 8'b00010010;
		color_arr[14988] = 8'b00010010;
		color_arr[14989] = 8'b00010010;
		color_arr[14990] = 8'b00010010;
		color_arr[14991] = 8'b00010010;
		color_arr[14992] = 8'b00010010;
		color_arr[14993] = 8'b00010010;
		color_arr[14994] = 8'b00100000;
		color_arr[14995] = 8'b00100000;
		color_arr[14996] = 8'b00100000;
		color_arr[14997] = 8'b00100000;
		color_arr[14998] = 8'b00100000;
		color_arr[14999] = 8'b00100000;
		color_arr[15000] = 8'b00100000;
		color_arr[15001] = 8'b00100000;
		color_arr[15002] = 8'b00100000;
		color_arr[15003] = 8'b00100000;
		color_arr[15004] = 8'b00100000;
		color_arr[15005] = 8'b00100000;
		color_arr[15006] = 8'b00100000;
		color_arr[15007] = 8'b00100000;
		color_arr[15008] = 8'b00100000;
		color_arr[15009] = 8'b00000000;
		color_arr[15010] = 8'b00000000;
		color_arr[15011] = 8'b00000000;
		color_arr[15012] = 8'b00000000;
		color_arr[15013] = 8'b00100000;
		color_arr[15014] = 8'b00100000;
		color_arr[15015] = 8'b00100000;
		color_arr[15016] = 8'b00100000;
		color_arr[15017] = 8'b00100000;
		color_arr[15018] = 8'b00100000;
		color_arr[15019] = 8'b00100000;
		color_arr[15020] = 8'b00100000;
		color_arr[15021] = 8'b00100000;
		color_arr[15022] = 8'b00100000;
		color_arr[15023] = 8'b00100000;
		color_arr[15024] = 8'b00100000;
		color_arr[15025] = 8'b00100000;
		color_arr[15026] = 8'b00100000;
		color_arr[15027] = 8'b00000000;
		color_arr[15028] = 8'b00000000;
		color_arr[15029] = 8'b00000000;
		color_arr[15030] = 8'b00000000;
		color_arr[15031] = 8'b00000000;
		color_arr[15032] = 8'b00100000;
		color_arr[15033] = 8'b00100000;
		color_arr[15034] = 8'b00100000;
		color_arr[15035] = 8'b00100000;
		color_arr[15036] = 8'b00100000;
		color_arr[15037] = 8'b00100000;
		color_arr[15038] = 8'b00100000;
		color_arr[15039] = 8'b00100000;
		color_arr[15040] = 8'b00100000;
		color_arr[15041] = 8'b00100000;
		color_arr[15042] = 8'b00100000;
		color_arr[15043] = 8'b00100000;
		color_arr[15044] = 8'b00100000;
		color_arr[15045] = 8'b00100000;
		color_arr[15046] = 8'b00100000;
		color_arr[15047] = 8'b00100000;
		color_arr[15048] = 8'b00100000;
		color_arr[15049] = 8'b00100000;
		color_arr[15050] = 8'b00100000;
		color_arr[15051] = 8'b00100000;
		color_arr[15052] = 8'b00100000;
		color_arr[15053] = 8'b00100000;
		color_arr[15054] = 8'b00100000;
		color_arr[15055] = 8'b00100000;
		color_arr[15056] = 8'b00100000;
		color_arr[15057] = 8'b00100000;
		color_arr[15058] = 8'b00100000;
		color_arr[15059] = 8'b00100000;
		color_arr[15060] = 8'b00100000;
		color_arr[15061] = 8'b00100000;
		color_arr[15062] = 8'b00100000;
		color_arr[15063] = 8'b00100000;
		color_arr[15064] = 8'b00100000;
		color_arr[15065] = 8'b00100000;
		color_arr[15066] = 8'b00100000;
		color_arr[15067] = 8'b00100000;
		color_arr[15068] = 8'b00100000;
		color_arr[15069] = 8'b00100000;
		color_arr[15070] = 8'b00100000;
		color_arr[15071] = 8'b00100000;
		color_arr[15072] = 8'b00100000;
		color_arr[15073] = 8'b00100000;
		color_arr[15074] = 8'b00100000;
		color_arr[15075] = 8'b00100000;
		color_arr[15076] = 8'b00100000;
		color_arr[15077] = 8'b00100000;
		color_arr[15078] = 8'b00100000;
		color_arr[15079] = 8'b00000000;
		color_arr[15080] = 8'b00000000;
		color_arr[15081] = 8'b00000000;
		color_arr[15082] = 8'b00000000;
		color_arr[15083] = 8'b00000000;
		color_arr[15084] = 8'b00000000;
		color_arr[15085] = 8'b00000000;
		color_arr[15086] = 8'b00100000;
		color_arr[15087] = 8'b00100000;
		color_arr[15088] = 8'b00100000;
		color_arr[15089] = 8'b00100000;
		color_arr[15090] = 8'b00100000;
		color_arr[15091] = 8'b00100000;
		color_arr[15092] = 8'b00100000;
		color_arr[15093] = 8'b00100000;
		color_arr[15094] = 8'b00100000;
		color_arr[15095] = 8'b00100000;
		color_arr[15096] = 8'b00100000;
		color_arr[15097] = 8'b00000000;
		color_arr[15098] = 8'b00000000;
		color_arr[15099] = 8'b00100000;
		color_arr[15100] = 8'b00100000;
		color_arr[15101] = 8'b00010010;
		color_arr[15102] = 8'b00010010;
		color_arr[15103] = 8'b00010010;
		color_arr[15104] = 8'b00010010;
		color_arr[15105] = 8'b00010010;
		color_arr[15106] = 8'b00010010;
		color_arr[15107] = 8'b00010010;
		color_arr[15108] = 8'b00000000;
		color_arr[15109] = 8'b00000000;
		color_arr[15110] = 8'b00000000;
		color_arr[15111] = 8'b00000000;
		color_arr[15112] = 8'b00000000;
		color_arr[15113] = 8'b00010010;
		color_arr[15114] = 8'b00010010;
		color_arr[15115] = 8'b00010010;
		color_arr[15116] = 8'b00010010;
		color_arr[15117] = 8'b00010010;
		color_arr[15118] = 8'b00010010;
		color_arr[15119] = 8'b00010010;
		color_arr[15120] = 8'b00010010;
		color_arr[15121] = 8'b00010010;
		color_arr[15122] = 8'b00100000;
		color_arr[15123] = 8'b00100000;
		color_arr[15124] = 8'b00100000;
		color_arr[15125] = 8'b00100000;
		color_arr[15126] = 8'b00100000;
		color_arr[15127] = 8'b00100000;
		color_arr[15128] = 8'b00100000;
		color_arr[15129] = 8'b00100000;
		color_arr[15130] = 8'b00100000;
		color_arr[15131] = 8'b00100000;
		color_arr[15132] = 8'b00100000;
		color_arr[15133] = 8'b00100000;
		color_arr[15134] = 8'b00100000;
		color_arr[15135] = 8'b00100000;
		color_arr[15136] = 8'b00000000;
		color_arr[15137] = 8'b00000000;
		color_arr[15138] = 8'b00000000;
		color_arr[15139] = 8'b00000000;
		color_arr[15140] = 8'b00100000;
		color_arr[15141] = 8'b00100000;
		color_arr[15142] = 8'b00100000;
		color_arr[15143] = 8'b00100000;
		color_arr[15144] = 8'b00100000;
		color_arr[15145] = 8'b00100000;
		color_arr[15146] = 8'b00100000;
		color_arr[15147] = 8'b00100000;
		color_arr[15148] = 8'b00100000;
		color_arr[15149] = 8'b00100000;
		color_arr[15150] = 8'b00100000;
		color_arr[15151] = 8'b00100000;
		color_arr[15152] = 8'b00100000;
		color_arr[15153] = 8'b00100000;
		color_arr[15154] = 8'b00000000;
		color_arr[15155] = 8'b00000000;
		color_arr[15156] = 8'b00000000;
		color_arr[15157] = 8'b00000000;
		color_arr[15158] = 8'b00100000;
		color_arr[15159] = 8'b00100000;
		color_arr[15160] = 8'b00100000;
		color_arr[15161] = 8'b00100000;
		color_arr[15162] = 8'b00100000;
		color_arr[15163] = 8'b00100000;
		color_arr[15164] = 8'b00100000;
		color_arr[15165] = 8'b00100000;
		color_arr[15166] = 8'b00100000;
		color_arr[15167] = 8'b00100000;
		color_arr[15168] = 8'b00100000;
		color_arr[15169] = 8'b00100000;
		color_arr[15170] = 8'b00100000;
		color_arr[15171] = 8'b00100000;
		color_arr[15172] = 8'b00100000;
		color_arr[15173] = 8'b00100000;
		color_arr[15174] = 8'b00100000;
		color_arr[15175] = 8'b00100000;
		color_arr[15176] = 8'b00100000;
		color_arr[15177] = 8'b00100000;
		color_arr[15178] = 8'b00100000;
		color_arr[15179] = 8'b00100000;
		color_arr[15180] = 8'b00100000;
		color_arr[15181] = 8'b00100000;
		color_arr[15182] = 8'b00100000;
		color_arr[15183] = 8'b00100000;
		color_arr[15184] = 8'b00100000;
		color_arr[15185] = 8'b00100000;
		color_arr[15186] = 8'b00100000;
		color_arr[15187] = 8'b00100000;
		color_arr[15188] = 8'b00100000;
		color_arr[15189] = 8'b00100000;
		color_arr[15190] = 8'b00100000;
		color_arr[15191] = 8'b00100000;
		color_arr[15192] = 8'b00100000;
		color_arr[15193] = 8'b00100000;
		color_arr[15194] = 8'b00100000;
		color_arr[15195] = 8'b00100000;
		color_arr[15196] = 8'b00100000;
		color_arr[15197] = 8'b00100000;
		color_arr[15198] = 8'b00100000;
		color_arr[15199] = 8'b00100000;
		color_arr[15200] = 8'b00100000;
		color_arr[15201] = 8'b00100000;
		color_arr[15202] = 8'b00100000;
		color_arr[15203] = 8'b00100000;
		color_arr[15204] = 8'b00100000;
		color_arr[15205] = 8'b00100000;
		color_arr[15206] = 8'b00100000;
		color_arr[15207] = 8'b00100000;
		color_arr[15208] = 8'b00100000;
		color_arr[15209] = 8'b00100000;
		color_arr[15210] = 8'b00000000;
		color_arr[15211] = 8'b00000000;
		color_arr[15212] = 8'b00000000;
		color_arr[15213] = 8'b00000000;
		color_arr[15214] = 8'b00000000;
		color_arr[15215] = 8'b00000000;
		color_arr[15216] = 8'b00000000;
		color_arr[15217] = 8'b00000000;
		color_arr[15218] = 8'b00100000;
		color_arr[15219] = 8'b00100000;
		color_arr[15220] = 8'b00100000;
		color_arr[15221] = 8'b00100000;
		color_arr[15222] = 8'b00100000;
		color_arr[15223] = 8'b00100000;
		color_arr[15224] = 8'b00100000;
		color_arr[15225] = 8'b00000000;
		color_arr[15226] = 8'b00000000;
		color_arr[15227] = 8'b00100000;
		color_arr[15228] = 8'b00100000;
		color_arr[15229] = 8'b00010010;
		color_arr[15230] = 8'b00010010;
		color_arr[15231] = 8'b00010010;
		color_arr[15232] = 8'b00010010;
		color_arr[15233] = 8'b00010010;
		color_arr[15234] = 8'b00010010;
		color_arr[15235] = 8'b00010010;
		color_arr[15236] = 8'b00010010;
		color_arr[15237] = 8'b00010010;
		color_arr[15238] = 8'b00000000;
		color_arr[15239] = 8'b00000000;
		color_arr[15240] = 8'b00000000;
		color_arr[15241] = 8'b00000000;
		color_arr[15242] = 8'b00000000;
		color_arr[15243] = 8'b00010010;
		color_arr[15244] = 8'b00010010;
		color_arr[15245] = 8'b00010010;
		color_arr[15246] = 8'b00010010;
		color_arr[15247] = 8'b00010010;
		color_arr[15248] = 8'b00010010;
		color_arr[15249] = 8'b00010010;
		color_arr[15250] = 8'b00100000;
		color_arr[15251] = 8'b00100000;
		color_arr[15252] = 8'b00100000;
		color_arr[15253] = 8'b00100000;
		color_arr[15254] = 8'b00100000;
		color_arr[15255] = 8'b00100000;
		color_arr[15256] = 8'b00100000;
		color_arr[15257] = 8'b00100000;
		color_arr[15258] = 8'b00100000;
		color_arr[15259] = 8'b00100000;
		color_arr[15260] = 8'b00100000;
		color_arr[15261] = 8'b00100000;
		color_arr[15262] = 8'b00100000;
		color_arr[15263] = 8'b00100000;
		color_arr[15264] = 8'b00000000;
		color_arr[15265] = 8'b00000000;
		color_arr[15266] = 8'b00100000;
		color_arr[15267] = 8'b00100000;
		color_arr[15268] = 8'b00100000;
		color_arr[15269] = 8'b00100000;
		color_arr[15270] = 8'b00100000;
		color_arr[15271] = 8'b00100000;
		color_arr[15272] = 8'b00100000;
		color_arr[15273] = 8'b00100000;
		color_arr[15274] = 8'b00100000;
		color_arr[15275] = 8'b00100000;
		color_arr[15276] = 8'b00100000;
		color_arr[15277] = 8'b00100000;
		color_arr[15278] = 8'b00100000;
		color_arr[15279] = 8'b00100000;
		color_arr[15280] = 8'b00000000;
		color_arr[15281] = 8'b00000000;
		color_arr[15282] = 8'b00000000;
		color_arr[15283] = 8'b00000000;
		color_arr[15284] = 8'b00100000;
		color_arr[15285] = 8'b00100000;
		color_arr[15286] = 8'b00100000;
		color_arr[15287] = 8'b00100000;
		color_arr[15288] = 8'b00100000;
		color_arr[15289] = 8'b00100000;
		color_arr[15290] = 8'b00100000;
		color_arr[15291] = 8'b00100000;
		color_arr[15292] = 8'b00100000;
		color_arr[15293] = 8'b00100000;
		color_arr[15294] = 8'b00100000;
		color_arr[15295] = 8'b00100000;
		color_arr[15296] = 8'b00100000;
		color_arr[15297] = 8'b00100000;
		color_arr[15298] = 8'b00100000;
		color_arr[15299] = 8'b00100000;
		color_arr[15300] = 8'b00100000;
		color_arr[15301] = 8'b00100000;
		color_arr[15302] = 8'b00100000;
		color_arr[15303] = 8'b00100000;
		color_arr[15304] = 8'b00100000;
		color_arr[15305] = 8'b00100000;
		color_arr[15306] = 8'b00100000;
		color_arr[15307] = 8'b00100000;
		color_arr[15308] = 8'b00100000;
		color_arr[15309] = 8'b00100000;
		color_arr[15310] = 8'b00100000;
		color_arr[15311] = 8'b00100000;
		color_arr[15312] = 8'b00100000;
		color_arr[15313] = 8'b00100000;
		color_arr[15314] = 8'b00100000;
		color_arr[15315] = 8'b00100000;
		color_arr[15316] = 8'b00100000;
		color_arr[15317] = 8'b00100000;
		color_arr[15318] = 8'b00100000;
		color_arr[15319] = 8'b00100000;
		color_arr[15320] = 8'b00100000;
		color_arr[15321] = 8'b00100000;
		color_arr[15322] = 8'b00100000;
		color_arr[15323] = 8'b00100000;
		color_arr[15324] = 8'b00100000;
		color_arr[15325] = 8'b00100000;
		color_arr[15326] = 8'b00100000;
		color_arr[15327] = 8'b00100000;
		color_arr[15328] = 8'b00100000;
		color_arr[15329] = 8'b00100000;
		color_arr[15330] = 8'b00100000;
		color_arr[15331] = 8'b00100000;
		color_arr[15332] = 8'b00100000;
		color_arr[15333] = 8'b00100000;
		color_arr[15334] = 8'b00100000;
		color_arr[15335] = 8'b00100000;
		color_arr[15336] = 8'b00100000;
		color_arr[15337] = 8'b00100000;
		color_arr[15338] = 8'b00100000;
		color_arr[15339] = 8'b00100000;
		color_arr[15340] = 8'b00100000;
		color_arr[15341] = 8'b00000000;
		color_arr[15342] = 8'b00000000;
		color_arr[15343] = 8'b00000000;
		color_arr[15344] = 8'b00000000;
		color_arr[15345] = 8'b00000000;
		color_arr[15346] = 8'b00000000;
		color_arr[15347] = 8'b00000000;
		color_arr[15348] = 8'b00000000;
		color_arr[15349] = 8'b00100000;
		color_arr[15350] = 8'b00100000;
		color_arr[15351] = 8'b00100000;
		color_arr[15352] = 8'b00100000;
		color_arr[15353] = 8'b00000000;
		color_arr[15354] = 8'b00000000;
		color_arr[15355] = 8'b00100000;
		color_arr[15356] = 8'b00100000;
		color_arr[15357] = 8'b00010010;
		color_arr[15358] = 8'b00010010;
		color_arr[15359] = 8'b00010010;
		color_arr[15360] = 8'b00010010;
		color_arr[15361] = 8'b00010010;
		color_arr[15362] = 8'b00010010;
		color_arr[15363] = 8'b00010010;
		color_arr[15364] = 8'b00010010;
		color_arr[15365] = 8'b00010010;
		color_arr[15366] = 8'b00010010;
		color_arr[15367] = 8'b00010010;
		color_arr[15368] = 8'b00000000;
		color_arr[15369] = 8'b00000000;
		color_arr[15370] = 8'b00000000;
		color_arr[15371] = 8'b00000000;
		color_arr[15372] = 8'b00000000;
		color_arr[15373] = 8'b00010010;
		color_arr[15374] = 8'b00010010;
		color_arr[15375] = 8'b00010010;
		color_arr[15376] = 8'b00010010;
		color_arr[15377] = 8'b00010010;
		color_arr[15378] = 8'b00100000;
		color_arr[15379] = 8'b00100000;
		color_arr[15380] = 8'b00100000;
		color_arr[15381] = 8'b00100000;
		color_arr[15382] = 8'b00100000;
		color_arr[15383] = 8'b00100000;
		color_arr[15384] = 8'b00100000;
		color_arr[15385] = 8'b00100000;
		color_arr[15386] = 8'b00100000;
		color_arr[15387] = 8'b00100000;
		color_arr[15388] = 8'b00100000;
		color_arr[15389] = 8'b00100000;
		color_arr[15390] = 8'b00100000;
		color_arr[15391] = 8'b00100000;
		color_arr[15392] = 8'b00100000;
		color_arr[15393] = 8'b00100000;
		color_arr[15394] = 8'b00100000;
		color_arr[15395] = 8'b00100000;
		color_arr[15396] = 8'b00100000;
		color_arr[15397] = 8'b00100000;
		color_arr[15398] = 8'b00100000;
		color_arr[15399] = 8'b00100000;
		color_arr[15400] = 8'b00100000;
		color_arr[15401] = 8'b00100000;
		color_arr[15402] = 8'b00100000;
		color_arr[15403] = 8'b00100000;
		color_arr[15404] = 8'b00100000;
		color_arr[15405] = 8'b00100000;
		color_arr[15406] = 8'b00100000;
		color_arr[15407] = 8'b00000000;
		color_arr[15408] = 8'b00000000;
		color_arr[15409] = 8'b00000000;
		color_arr[15410] = 8'b00000000;
		color_arr[15411] = 8'b00100000;
		color_arr[15412] = 8'b00100000;
		color_arr[15413] = 8'b00100000;
		color_arr[15414] = 8'b00100000;
		color_arr[15415] = 8'b00100000;
		color_arr[15416] = 8'b00100000;
		color_arr[15417] = 8'b00100000;
		color_arr[15418] = 8'b00100000;
		color_arr[15419] = 8'b00100000;
		color_arr[15420] = 8'b00100000;
		color_arr[15421] = 8'b00100000;
		color_arr[15422] = 8'b00100000;
		color_arr[15423] = 8'b00100000;
		color_arr[15424] = 8'b00100000;
		color_arr[15425] = 8'b00100000;
		color_arr[15426] = 8'b00100000;
		color_arr[15427] = 8'b00100000;
		color_arr[15428] = 8'b00100000;
		color_arr[15429] = 8'b00100000;
		color_arr[15430] = 8'b00100000;
		color_arr[15431] = 8'b00100000;
		color_arr[15432] = 8'b00100000;
		color_arr[15433] = 8'b00100000;
		color_arr[15434] = 8'b00100000;
		color_arr[15435] = 8'b00100000;
		color_arr[15436] = 8'b00100000;
		color_arr[15437] = 8'b00100000;
		color_arr[15438] = 8'b00100000;
		color_arr[15439] = 8'b00100000;
		color_arr[15440] = 8'b00100000;
		color_arr[15441] = 8'b00100000;
		color_arr[15442] = 8'b00100000;
		color_arr[15443] = 8'b00100000;
		color_arr[15444] = 8'b00100000;
		color_arr[15445] = 8'b00100000;
		color_arr[15446] = 8'b00100000;
		color_arr[15447] = 8'b00100000;
		color_arr[15448] = 8'b00100000;
		color_arr[15449] = 8'b00100000;
		color_arr[15450] = 8'b00100000;
		color_arr[15451] = 8'b00100000;
		color_arr[15452] = 8'b00100000;
		color_arr[15453] = 8'b00100000;
		color_arr[15454] = 8'b00100000;
		color_arr[15455] = 8'b00100000;
		color_arr[15456] = 8'b00100000;
		color_arr[15457] = 8'b00100000;
		color_arr[15458] = 8'b00100000;
		color_arr[15459] = 8'b00100000;
		color_arr[15460] = 8'b00100000;
		color_arr[15461] = 8'b00100000;
		color_arr[15462] = 8'b00100000;
		color_arr[15463] = 8'b00100000;
		color_arr[15464] = 8'b00100000;
		color_arr[15465] = 8'b00100000;
		color_arr[15466] = 8'b00100000;
		color_arr[15467] = 8'b00100000;
		color_arr[15468] = 8'b00100000;
		color_arr[15469] = 8'b00100000;
		color_arr[15470] = 8'b00100000;
		color_arr[15471] = 8'b00100000;
		color_arr[15472] = 8'b00100000;
		color_arr[15473] = 8'b00000000;
		color_arr[15474] = 8'b00000000;
		color_arr[15475] = 8'b00000000;
		color_arr[15476] = 8'b00000000;
		color_arr[15477] = 8'b00000000;
		color_arr[15478] = 8'b00000000;
		color_arr[15479] = 8'b00000000;
		color_arr[15480] = 8'b00100000;
		color_arr[15481] = 8'b00000000;
		color_arr[15482] = 8'b00000000;
		color_arr[15483] = 8'b00100000;
		color_arr[15484] = 8'b00100000;
		color_arr[15485] = 8'b00010010;
		color_arr[15486] = 8'b00010010;
		color_arr[15487] = 8'b00010010;
		color_arr[15488] = 8'b00010010;
		color_arr[15489] = 8'b00010010;
		color_arr[15490] = 8'b00010010;
		color_arr[15491] = 8'b00010010;
		color_arr[15492] = 8'b00010010;
		color_arr[15493] = 8'b00010010;
		color_arr[15494] = 8'b00010010;
		color_arr[15495] = 8'b00010010;
		color_arr[15496] = 8'b00010010;
		color_arr[15497] = 8'b00010010;
		color_arr[15498] = 8'b00000000;
		color_arr[15499] = 8'b00000000;
		color_arr[15500] = 8'b00000000;
		color_arr[15501] = 8'b00000000;
		color_arr[15502] = 8'b00000000;
		color_arr[15503] = 8'b00000000;
		color_arr[15504] = 8'b00010010;
		color_arr[15505] = 8'b00010010;
		color_arr[15506] = 8'b00010010;
		color_arr[15507] = 8'b00010010;
		color_arr[15508] = 8'b00010010;
		color_arr[15509] = 8'b00010010;
		color_arr[15510] = 8'b00010010;
		color_arr[15511] = 8'b00010010;
		color_arr[15512] = 8'b00010010;
		color_arr[15513] = 8'b00010010;
		color_arr[15514] = 8'b00010010;
		color_arr[15515] = 8'b00010010;
		color_arr[15516] = 8'b00010010;
		color_arr[15517] = 8'b00010010;
		color_arr[15518] = 8'b00010010;
		color_arr[15519] = 8'b00010010;
		color_arr[15520] = 8'b00010010;
		color_arr[15521] = 8'b00010010;
		color_arr[15522] = 8'b00010010;
		color_arr[15523] = 8'b00010010;
		color_arr[15524] = 8'b00010010;
		color_arr[15525] = 8'b00010010;
		color_arr[15526] = 8'b00010010;
		color_arr[15527] = 8'b00010010;
		color_arr[15528] = 8'b00010010;
		color_arr[15529] = 8'b00010010;
		color_arr[15530] = 8'b00010010;
		color_arr[15531] = 8'b00010010;
		color_arr[15532] = 8'b00010010;
		color_arr[15533] = 8'b00000000;
		color_arr[15534] = 8'b00000000;
		color_arr[15535] = 8'b00000000;
		color_arr[15536] = 8'b00000000;
		color_arr[15537] = 8'b00010010;
		color_arr[15538] = 8'b00010010;
		color_arr[15539] = 8'b00010010;
		color_arr[15540] = 8'b00010010;
		color_arr[15541] = 8'b00010010;
		color_arr[15542] = 8'b00010010;
		color_arr[15543] = 8'b00010010;
		color_arr[15544] = 8'b00010010;
		color_arr[15545] = 8'b00010010;
		color_arr[15546] = 8'b00010010;
		color_arr[15547] = 8'b00010010;
		color_arr[15548] = 8'b00010010;
		color_arr[15549] = 8'b00010010;
		color_arr[15550] = 8'b00010010;
		color_arr[15551] = 8'b00010010;
		color_arr[15552] = 8'b00010010;
		color_arr[15553] = 8'b00010010;
		color_arr[15554] = 8'b00010010;
		color_arr[15555] = 8'b00010010;
		color_arr[15556] = 8'b00010010;
		color_arr[15557] = 8'b00010010;
		color_arr[15558] = 8'b00010010;
		color_arr[15559] = 8'b00010010;
		color_arr[15560] = 8'b00010010;
		color_arr[15561] = 8'b00010010;
		color_arr[15562] = 8'b00010010;
		color_arr[15563] = 8'b00010010;
		color_arr[15564] = 8'b00010010;
		color_arr[15565] = 8'b00010010;
		color_arr[15566] = 8'b00010010;
		color_arr[15567] = 8'b00010010;
		color_arr[15568] = 8'b00010010;
		color_arr[15569] = 8'b00010010;
		color_arr[15570] = 8'b00010010;
		color_arr[15571] = 8'b00010010;
		color_arr[15572] = 8'b00010010;
		color_arr[15573] = 8'b00010010;
		color_arr[15574] = 8'b00010010;
		color_arr[15575] = 8'b00010010;
		color_arr[15576] = 8'b00010010;
		color_arr[15577] = 8'b00010010;
		color_arr[15578] = 8'b00010010;
		color_arr[15579] = 8'b00010010;
		color_arr[15580] = 8'b00010010;
		color_arr[15581] = 8'b00010010;
		color_arr[15582] = 8'b00010010;
		color_arr[15583] = 8'b00010010;
		color_arr[15584] = 8'b00010010;
		color_arr[15585] = 8'b00010010;
		color_arr[15586] = 8'b00010010;
		color_arr[15587] = 8'b00010010;
		color_arr[15588] = 8'b00010010;
		color_arr[15589] = 8'b00010010;
		color_arr[15590] = 8'b00010010;
		color_arr[15591] = 8'b00010010;
		color_arr[15592] = 8'b00010010;
		color_arr[15593] = 8'b00010010;
		color_arr[15594] = 8'b00010010;
		color_arr[15595] = 8'b00010010;
		color_arr[15596] = 8'b00010010;
		color_arr[15597] = 8'b00010010;
		color_arr[15598] = 8'b00010010;
		color_arr[15599] = 8'b00010010;
		color_arr[15600] = 8'b00010010;
		color_arr[15601] = 8'b00010010;
		color_arr[15602] = 8'b00010010;
		color_arr[15603] = 8'b00010010;
		color_arr[15604] = 8'b00000000;
		color_arr[15605] = 8'b00000000;
		color_arr[15606] = 8'b00000000;
		color_arr[15607] = 8'b00000000;
		color_arr[15608] = 8'b00000000;
		color_arr[15609] = 8'b00000000;
		color_arr[15610] = 8'b00000000;
		color_arr[15611] = 8'b00010010;
		color_arr[15612] = 8'b00010010;
		color_arr[15613] = 8'b00010010;
		color_arr[15614] = 8'b00010010;
		color_arr[15615] = 8'b00010010;
		color_arr[15616] = 8'b00010010;
		color_arr[15617] = 8'b00010010;
		color_arr[15618] = 8'b00010010;
		color_arr[15619] = 8'b00010010;
		color_arr[15620] = 8'b00010010;
		color_arr[15621] = 8'b00010010;
		color_arr[15622] = 8'b00010010;
		color_arr[15623] = 8'b00010010;
		color_arr[15624] = 8'b00010010;
		color_arr[15625] = 8'b00010010;
		color_arr[15626] = 8'b00010010;
		color_arr[15627] = 8'b00010010;
		color_arr[15628] = 8'b00000000;
		color_arr[15629] = 8'b00000000;
		color_arr[15630] = 8'b00000000;
		color_arr[15631] = 8'b00000000;
		color_arr[15632] = 8'b00000000;
		color_arr[15633] = 8'b00000000;
		color_arr[15634] = 8'b00010010;
		color_arr[15635] = 8'b00010010;
		color_arr[15636] = 8'b00010010;
		color_arr[15637] = 8'b00010010;
		color_arr[15638] = 8'b00010010;
		color_arr[15639] = 8'b00010010;
		color_arr[15640] = 8'b00010010;
		color_arr[15641] = 8'b00010010;
		color_arr[15642] = 8'b00010010;
		color_arr[15643] = 8'b00010010;
		color_arr[15644] = 8'b00010010;
		color_arr[15645] = 8'b00010010;
		color_arr[15646] = 8'b00010010;
		color_arr[15647] = 8'b00010010;
		color_arr[15648] = 8'b00010010;
		color_arr[15649] = 8'b00010010;
		color_arr[15650] = 8'b00010010;
		color_arr[15651] = 8'b00010010;
		color_arr[15652] = 8'b00010010;
		color_arr[15653] = 8'b00010010;
		color_arr[15654] = 8'b00010010;
		color_arr[15655] = 8'b00010010;
		color_arr[15656] = 8'b00010010;
		color_arr[15657] = 8'b00010010;
		color_arr[15658] = 8'b00010010;
		color_arr[15659] = 8'b00010010;
		color_arr[15660] = 8'b00000000;
		color_arr[15661] = 8'b00000000;
		color_arr[15662] = 8'b00000000;
		color_arr[15663] = 8'b00000000;
		color_arr[15664] = 8'b00010010;
		color_arr[15665] = 8'b00010010;
		color_arr[15666] = 8'b00010010;
		color_arr[15667] = 8'b00010010;
		color_arr[15668] = 8'b00010010;
		color_arr[15669] = 8'b00010010;
		color_arr[15670] = 8'b00010010;
		color_arr[15671] = 8'b00010010;
		color_arr[15672] = 8'b00010010;
		color_arr[15673] = 8'b00010010;
		color_arr[15674] = 8'b00010010;
		color_arr[15675] = 8'b00010010;
		color_arr[15676] = 8'b00010010;
		color_arr[15677] = 8'b00010010;
		color_arr[15678] = 8'b00010010;
		color_arr[15679] = 8'b00010010;
		color_arr[15680] = 8'b00010010;
		color_arr[15681] = 8'b00010010;
		color_arr[15682] = 8'b00010010;
		color_arr[15683] = 8'b00010010;
		color_arr[15684] = 8'b00010010;
		color_arr[15685] = 8'b00010010;
		color_arr[15686] = 8'b00010010;
		color_arr[15687] = 8'b00010010;
		color_arr[15688] = 8'b00010010;
		color_arr[15689] = 8'b00010010;
		color_arr[15690] = 8'b00010010;
		color_arr[15691] = 8'b00010010;
		color_arr[15692] = 8'b00010010;
		color_arr[15693] = 8'b00010010;
		color_arr[15694] = 8'b00010010;
		color_arr[15695] = 8'b00010010;
		color_arr[15696] = 8'b00010010;
		color_arr[15697] = 8'b00010010;
		color_arr[15698] = 8'b00010010;
		color_arr[15699] = 8'b00010010;
		color_arr[15700] = 8'b00010010;
		color_arr[15701] = 8'b00010010;
		color_arr[15702] = 8'b00010010;
		color_arr[15703] = 8'b00010010;
		color_arr[15704] = 8'b00010010;
		color_arr[15705] = 8'b00010010;
		color_arr[15706] = 8'b00010010;
		color_arr[15707] = 8'b00010010;
		color_arr[15708] = 8'b00010010;
		color_arr[15709] = 8'b00010010;
		color_arr[15710] = 8'b00010010;
		color_arr[15711] = 8'b00010010;
		color_arr[15712] = 8'b00010010;
		color_arr[15713] = 8'b00010010;
		color_arr[15714] = 8'b00010010;
		color_arr[15715] = 8'b00010010;
		color_arr[15716] = 8'b00010010;
		color_arr[15717] = 8'b00010010;
		color_arr[15718] = 8'b00010010;
		color_arr[15719] = 8'b00010010;
		color_arr[15720] = 8'b00010010;
		color_arr[15721] = 8'b00010010;
		color_arr[15722] = 8'b00010010;
		color_arr[15723] = 8'b00010010;
		color_arr[15724] = 8'b00010010;
		color_arr[15725] = 8'b00010010;
		color_arr[15726] = 8'b00010010;
		color_arr[15727] = 8'b00010010;
		color_arr[15728] = 8'b00010010;
		color_arr[15729] = 8'b00010010;
		color_arr[15730] = 8'b00010010;
		color_arr[15731] = 8'b00010010;
		color_arr[15732] = 8'b00010010;
		color_arr[15733] = 8'b00010010;
		color_arr[15734] = 8'b00010010;
		color_arr[15735] = 8'b00000000;
		color_arr[15736] = 8'b00000000;
		color_arr[15737] = 8'b00000000;
		color_arr[15738] = 8'b00000000;
		color_arr[15739] = 8'b00010010;
		color_arr[15740] = 8'b00010010;
		color_arr[15741] = 8'b00010010;
		color_arr[15742] = 8'b00010010;
		color_arr[15743] = 8'b00010010;
		color_arr[15744] = 8'b00010010;
		color_arr[15745] = 8'b00010010;
		color_arr[15746] = 8'b00010010;
		color_arr[15747] = 8'b00010010;
		color_arr[15748] = 8'b00010010;
		color_arr[15749] = 8'b00010010;
		color_arr[15750] = 8'b00010010;
		color_arr[15751] = 8'b00010010;
		color_arr[15752] = 8'b00010010;
		color_arr[15753] = 8'b00010010;
		color_arr[15754] = 8'b00010010;
		color_arr[15755] = 8'b00010010;
		color_arr[15756] = 8'b00010010;
		color_arr[15757] = 8'b00010010;
		color_arr[15758] = 8'b00010010;
		color_arr[15759] = 8'b00000000;
		color_arr[15760] = 8'b00000000;
		color_arr[15761] = 8'b00000000;
		color_arr[15762] = 8'b00000000;
		color_arr[15763] = 8'b00000000;
		color_arr[15764] = 8'b00000000;
		color_arr[15765] = 8'b00010010;
		color_arr[15766] = 8'b00010010;
		color_arr[15767] = 8'b00010010;
		color_arr[15768] = 8'b00010010;
		color_arr[15769] = 8'b00010010;
		color_arr[15770] = 8'b00010010;
		color_arr[15771] = 8'b00010010;
		color_arr[15772] = 8'b00010010;
		color_arr[15773] = 8'b00010010;
		color_arr[15774] = 8'b00010010;
		color_arr[15775] = 8'b00010010;
		color_arr[15776] = 8'b00010010;
		color_arr[15777] = 8'b00010010;
		color_arr[15778] = 8'b00010010;
		color_arr[15779] = 8'b00010010;
		color_arr[15780] = 8'b00010010;
		color_arr[15781] = 8'b00010010;
		color_arr[15782] = 8'b00010010;
		color_arr[15783] = 8'b00010010;
		color_arr[15784] = 8'b00010010;
		color_arr[15785] = 8'b00010010;
		color_arr[15786] = 8'b00000000;
		color_arr[15787] = 8'b00000000;
		color_arr[15788] = 8'b00000000;
		color_arr[15789] = 8'b00000000;
		color_arr[15790] = 8'b00010010;
		color_arr[15791] = 8'b00010010;
		color_arr[15792] = 8'b00010010;
		color_arr[15793] = 8'b00010010;
		color_arr[15794] = 8'b00010010;
		color_arr[15795] = 8'b00010010;
		color_arr[15796] = 8'b00010010;
		color_arr[15797] = 8'b00010010;
		color_arr[15798] = 8'b00010010;
		color_arr[15799] = 8'b00010010;
		color_arr[15800] = 8'b00010010;
		color_arr[15801] = 8'b00010010;
		color_arr[15802] = 8'b00010010;
		color_arr[15803] = 8'b00010010;
		color_arr[15804] = 8'b00010010;
		color_arr[15805] = 8'b00010010;
		color_arr[15806] = 8'b00010010;
		color_arr[15807] = 8'b00010010;
		color_arr[15808] = 8'b00010010;
		color_arr[15809] = 8'b00010010;
		color_arr[15810] = 8'b00010010;
		color_arr[15811] = 8'b00010010;
		color_arr[15812] = 8'b00010010;
		color_arr[15813] = 8'b00010010;
		color_arr[15814] = 8'b00010010;
		color_arr[15815] = 8'b00010010;
		color_arr[15816] = 8'b00010010;
		color_arr[15817] = 8'b00010010;
		color_arr[15818] = 8'b00010010;
		color_arr[15819] = 8'b00010010;
		color_arr[15820] = 8'b00010010;
		color_arr[15821] = 8'b00010010;
		color_arr[15822] = 8'b00010010;
		color_arr[15823] = 8'b00010010;
		color_arr[15824] = 8'b00010010;
		color_arr[15825] = 8'b00010010;
		color_arr[15826] = 8'b00010010;
		color_arr[15827] = 8'b00010010;
		color_arr[15828] = 8'b00010010;
		color_arr[15829] = 8'b00010010;
		color_arr[15830] = 8'b00010010;
		color_arr[15831] = 8'b00010010;
		color_arr[15832] = 8'b00010010;
		color_arr[15833] = 8'b00010010;
		color_arr[15834] = 8'b00010010;
		color_arr[15835] = 8'b00010010;
		color_arr[15836] = 8'b00010010;
		color_arr[15837] = 8'b00010010;
		color_arr[15838] = 8'b00010010;
		color_arr[15839] = 8'b00010010;
		color_arr[15840] = 8'b00010010;
		color_arr[15841] = 8'b00010010;
		color_arr[15842] = 8'b00010010;
		color_arr[15843] = 8'b00010010;
		color_arr[15844] = 8'b00010010;
		color_arr[15845] = 8'b00010010;
		color_arr[15846] = 8'b00010010;
		color_arr[15847] = 8'b00010010;
		color_arr[15848] = 8'b00010010;
		color_arr[15849] = 8'b00010010;
		color_arr[15850] = 8'b00010010;
		color_arr[15851] = 8'b00010010;
		color_arr[15852] = 8'b00010010;
		color_arr[15853] = 8'b00010010;
		color_arr[15854] = 8'b00010010;
		color_arr[15855] = 8'b00010010;
		color_arr[15856] = 8'b00010010;
		color_arr[15857] = 8'b00010010;
		color_arr[15858] = 8'b00010010;
		color_arr[15859] = 8'b00010010;
		color_arr[15860] = 8'b00010010;
		color_arr[15861] = 8'b00010010;
		color_arr[15862] = 8'b00010010;
		color_arr[15863] = 8'b00010010;
		color_arr[15864] = 8'b00010010;
		color_arr[15865] = 8'b00010010;
		color_arr[15866] = 8'b00010010;
		color_arr[15867] = 8'b00010010;
		color_arr[15868] = 8'b00010010;
		color_arr[15869] = 8'b00010010;
		color_arr[15870] = 8'b00010010;
		color_arr[15871] = 8'b00010010;
		color_arr[15872] = 8'b00010010;
		color_arr[15873] = 8'b00010010;
		color_arr[15874] = 8'b00010010;
		color_arr[15875] = 8'b00010010;
		color_arr[15876] = 8'b00010010;
		color_arr[15877] = 8'b00010010;
		color_arr[15878] = 8'b00010010;
		color_arr[15879] = 8'b00010010;
		color_arr[15880] = 8'b00010010;
		color_arr[15881] = 8'b00010010;
		color_arr[15882] = 8'b00010010;
		color_arr[15883] = 8'b00010010;
		color_arr[15884] = 8'b00010010;
		color_arr[15885] = 8'b00010010;
		color_arr[15886] = 8'b00010010;
		color_arr[15887] = 8'b00010010;
		color_arr[15888] = 8'b00010010;
		color_arr[15889] = 8'b00000000;
		color_arr[15890] = 8'b00000000;
		color_arr[15891] = 8'b00000000;
		color_arr[15892] = 8'b00000000;
		color_arr[15893] = 8'b00000000;
		color_arr[15894] = 8'b00000000;
		color_arr[15895] = 8'b00000000;
		color_arr[15896] = 8'b00010010;
		color_arr[15897] = 8'b00010010;
		color_arr[15898] = 8'b00010010;
		color_arr[15899] = 8'b00010010;
		color_arr[15900] = 8'b00010010;
		color_arr[15901] = 8'b00010010;
		color_arr[15902] = 8'b00010010;
		color_arr[15903] = 8'b00010010;
		color_arr[15904] = 8'b00010010;
		color_arr[15905] = 8'b00010010;
		color_arr[15906] = 8'b00010010;
		color_arr[15907] = 8'b00010010;
		color_arr[15908] = 8'b00010010;
		color_arr[15909] = 8'b00010010;
		color_arr[15910] = 8'b00010010;
		color_arr[15911] = 8'b00010010;
		color_arr[15912] = 8'b00010010;
		color_arr[15913] = 8'b00000000;
		color_arr[15914] = 8'b00000000;
		color_arr[15915] = 8'b00000000;
		color_arr[15916] = 8'b00000000;
		color_arr[15917] = 8'b00010010;
		color_arr[15918] = 8'b00010010;
		color_arr[15919] = 8'b00010010;
		color_arr[15920] = 8'b00010010;
		color_arr[15921] = 8'b00010010;
		color_arr[15922] = 8'b00010010;
		color_arr[15923] = 8'b00010010;
		color_arr[15924] = 8'b00010010;
		color_arr[15925] = 8'b00010010;
		color_arr[15926] = 8'b00010010;
		color_arr[15927] = 8'b00010010;
		color_arr[15928] = 8'b00010010;
		color_arr[15929] = 8'b00010010;
		color_arr[15930] = 8'b00010010;
		color_arr[15931] = 8'b00010010;
		color_arr[15932] = 8'b00010010;
		color_arr[15933] = 8'b00010010;
		color_arr[15934] = 8'b00010010;
		color_arr[15935] = 8'b00010010;
		color_arr[15936] = 8'b00010010;
		color_arr[15937] = 8'b00010010;
		color_arr[15938] = 8'b00010010;
		color_arr[15939] = 8'b00010010;
		color_arr[15940] = 8'b00010010;
		color_arr[15941] = 8'b00010010;
		color_arr[15942] = 8'b00010010;
		color_arr[15943] = 8'b00010010;
		color_arr[15944] = 8'b00010010;
		color_arr[15945] = 8'b00010010;
		color_arr[15946] = 8'b00010010;
		color_arr[15947] = 8'b00010010;
		color_arr[15948] = 8'b00010010;
		color_arr[15949] = 8'b00010010;
		color_arr[15950] = 8'b00010010;
		color_arr[15951] = 8'b00010010;
		color_arr[15952] = 8'b00010010;
		color_arr[15953] = 8'b00010010;
		color_arr[15954] = 8'b00010010;
		color_arr[15955] = 8'b00010010;
		color_arr[15956] = 8'b00010010;
		color_arr[15957] = 8'b00010010;
		color_arr[15958] = 8'b00010010;
		color_arr[15959] = 8'b00010010;
		color_arr[15960] = 8'b00010010;
		color_arr[15961] = 8'b00010010;
		color_arr[15962] = 8'b00010010;
		color_arr[15963] = 8'b00010010;
		color_arr[15964] = 8'b00010010;
		color_arr[15965] = 8'b00010010;
		color_arr[15966] = 8'b00010010;
		color_arr[15967] = 8'b00010010;
		color_arr[15968] = 8'b00010010;
		color_arr[15969] = 8'b00010010;
		color_arr[15970] = 8'b00010010;
		color_arr[15971] = 8'b00010010;
		color_arr[15972] = 8'b00010010;
		color_arr[15973] = 8'b00010010;
		color_arr[15974] = 8'b00010010;
		color_arr[15975] = 8'b00010010;
		color_arr[15976] = 8'b00010010;
		color_arr[15977] = 8'b00010010;
		color_arr[15978] = 8'b00010010;
		color_arr[15979] = 8'b00010010;
		color_arr[15980] = 8'b00010010;
		color_arr[15981] = 8'b00010010;
		color_arr[15982] = 8'b00010010;
		color_arr[15983] = 8'b00010010;
		color_arr[15984] = 8'b00010010;
		color_arr[15985] = 8'b00010010;
		color_arr[15986] = 8'b00010010;
		color_arr[15987] = 8'b00010010;
		color_arr[15988] = 8'b00010010;
		color_arr[15989] = 8'b00010010;
		color_arr[15990] = 8'b00010010;
		color_arr[15991] = 8'b00010010;
		color_arr[15992] = 8'b00010010;
		color_arr[15993] = 8'b00010010;
		color_arr[15994] = 8'b00010010;
		color_arr[15995] = 8'b00010010;
		color_arr[15996] = 8'b00010010;
		color_arr[15997] = 8'b00010010;
		color_arr[15998] = 8'b00010010;
		color_arr[15999] = 8'b00010010;
		color_arr[16000] = 8'b00010010;
		color_arr[16001] = 8'b00010010;
		color_arr[16002] = 8'b00010010;
		color_arr[16003] = 8'b00010010;
		color_arr[16004] = 8'b00010010;
		color_arr[16005] = 8'b00010010;
		color_arr[16006] = 8'b00010010;
		color_arr[16007] = 8'b00010010;
		color_arr[16008] = 8'b00010010;
		color_arr[16009] = 8'b00010010;
		color_arr[16010] = 8'b00010010;
		color_arr[16011] = 8'b00010010;
		color_arr[16012] = 8'b00010010;
		color_arr[16013] = 8'b00010010;
		color_arr[16014] = 8'b00010010;
		color_arr[16015] = 8'b00010010;
		color_arr[16016] = 8'b00010010;
		color_arr[16017] = 8'b00010010;
		color_arr[16018] = 8'b00010010;
		color_arr[16019] = 8'b00010010;
		color_arr[16020] = 8'b00000000;
		color_arr[16021] = 8'b00000000;
		color_arr[16022] = 8'b00000000;
		color_arr[16023] = 8'b00000000;
		color_arr[16024] = 8'b00010010;
		color_arr[16025] = 8'b00010010;
		color_arr[16026] = 8'b00010010;
		color_arr[16027] = 8'b00010010;
		color_arr[16028] = 8'b00010010;
		color_arr[16029] = 8'b00010010;
		color_arr[16030] = 8'b00010010;
		color_arr[16031] = 8'b00010010;
		color_arr[16032] = 8'b00010010;
		color_arr[16033] = 8'b00010010;
		color_arr[16034] = 8'b00010010;
		color_arr[16035] = 8'b00010010;
		color_arr[16036] = 8'b00010010;
		color_arr[16037] = 8'b00010010;
		color_arr[16038] = 8'b00010010;
		color_arr[16039] = 8'b00000000;
		color_arr[16040] = 8'b00000000;
		color_arr[16041] = 8'b00000000;
		color_arr[16042] = 8'b00000000;
		color_arr[16043] = 8'b00010010;
		color_arr[16044] = 8'b00010010;
		color_arr[16045] = 8'b00010010;
		color_arr[16046] = 8'b00010010;
		color_arr[16047] = 8'b00010010;
		color_arr[16048] = 8'b00010010;
		color_arr[16049] = 8'b00010010;
		color_arr[16050] = 8'b00010010;
		color_arr[16051] = 8'b00010010;
		color_arr[16052] = 8'b00010010;
		color_arr[16053] = 8'b00010010;
		color_arr[16054] = 8'b00010010;
		color_arr[16055] = 8'b00010010;
		color_arr[16056] = 8'b00010010;
		color_arr[16057] = 8'b00010010;
		color_arr[16058] = 8'b00010010;
		color_arr[16059] = 8'b00010010;
		color_arr[16060] = 8'b00010010;
		color_arr[16061] = 8'b00010010;
		color_arr[16062] = 8'b00010010;
		color_arr[16063] = 8'b00010010;
		color_arr[16064] = 8'b00010010;
		color_arr[16065] = 8'b00010010;
		color_arr[16066] = 8'b00010010;
		color_arr[16067] = 8'b00010010;
		color_arr[16068] = 8'b00010010;
		color_arr[16069] = 8'b00010010;
		color_arr[16070] = 8'b00010010;
		color_arr[16071] = 8'b00010010;
		color_arr[16072] = 8'b00010010;
		color_arr[16073] = 8'b00010010;
		color_arr[16074] = 8'b00010010;
		color_arr[16075] = 8'b00010010;
		color_arr[16076] = 8'b00010010;
		color_arr[16077] = 8'b00010010;
		color_arr[16078] = 8'b00010010;
		color_arr[16079] = 8'b00010010;
		color_arr[16080] = 8'b00010010;
		color_arr[16081] = 8'b00010010;
		color_arr[16082] = 8'b00010010;
		color_arr[16083] = 8'b00010010;
		color_arr[16084] = 8'b00010010;
		color_arr[16085] = 8'b00010010;
		color_arr[16086] = 8'b00010010;
		color_arr[16087] = 8'b00010010;
		color_arr[16088] = 8'b00010010;
		color_arr[16089] = 8'b00010010;
		color_arr[16090] = 8'b00010010;
		color_arr[16091] = 8'b00010010;
		color_arr[16092] = 8'b00010010;
		color_arr[16093] = 8'b00010010;
		color_arr[16094] = 8'b00010010;
		color_arr[16095] = 8'b00010010;
		color_arr[16096] = 8'b00010010;
		color_arr[16097] = 8'b00010010;
		color_arr[16098] = 8'b00010010;
		color_arr[16099] = 8'b00010010;
		color_arr[16100] = 8'b00010010;
		color_arr[16101] = 8'b00010010;
		color_arr[16102] = 8'b00010010;
		color_arr[16103] = 8'b00010010;
		color_arr[16104] = 8'b00010010;
		color_arr[16105] = 8'b00010010;
		color_arr[16106] = 8'b00010010;
		color_arr[16107] = 8'b00010010;
		color_arr[16108] = 8'b00010010;
		color_arr[16109] = 8'b00010010;
		color_arr[16110] = 8'b00010010;
		color_arr[16111] = 8'b00010010;
		color_arr[16112] = 8'b00010010;
		color_arr[16113] = 8'b00010010;
		color_arr[16114] = 8'b00010010;
		color_arr[16115] = 8'b00010010;
		color_arr[16116] = 8'b00010010;
		color_arr[16117] = 8'b00010010;
		color_arr[16118] = 8'b00010010;
		color_arr[16119] = 8'b00010010;
		color_arr[16120] = 8'b00010010;
		color_arr[16121] = 8'b00010010;
		color_arr[16122] = 8'b00010010;
		color_arr[16123] = 8'b00010010;
		color_arr[16124] = 8'b00010010;
		color_arr[16125] = 8'b00010010;
		color_arr[16126] = 8'b00010010;
		color_arr[16127] = 8'b00010010;
		color_arr[16128] = 8'b00010010;
		color_arr[16129] = 8'b00010010;
		color_arr[16130] = 8'b00010010;
		color_arr[16131] = 8'b00010010;
		color_arr[16132] = 8'b00010010;
		color_arr[16133] = 8'b00010010;
		color_arr[16134] = 8'b00010010;
		color_arr[16135] = 8'b00010010;
		color_arr[16136] = 8'b00010010;
		color_arr[16137] = 8'b00010010;
		color_arr[16138] = 8'b00010010;
		color_arr[16139] = 8'b00010010;
		color_arr[16140] = 8'b00010010;
		color_arr[16141] = 8'b00010010;
		color_arr[16142] = 8'b00010010;
		color_arr[16143] = 8'b00010010;
		color_arr[16144] = 8'b00010010;
		color_arr[16145] = 8'b00010010;
		color_arr[16146] = 8'b00010010;
		color_arr[16147] = 8'b00010010;
		color_arr[16148] = 8'b00010010;
		color_arr[16149] = 8'b00010010;
		color_arr[16150] = 8'b00000000;
		color_arr[16151] = 8'b00000000;
		color_arr[16152] = 8'b00010010;
		color_arr[16153] = 8'b00010010;
		color_arr[16154] = 8'b00010010;
		color_arr[16155] = 8'b00010010;
		color_arr[16156] = 8'b00010010;
		color_arr[16157] = 8'b00010010;
		color_arr[16158] = 8'b00010010;
		color_arr[16159] = 8'b00010010;
		color_arr[16160] = 8'b00010010;
		color_arr[16161] = 8'b00010010;
		color_arr[16162] = 8'b00010010;
		color_arr[16163] = 8'b00010010;
		color_arr[16164] = 8'b00010010;
		color_arr[16165] = 8'b00000000;
		color_arr[16166] = 8'b00000000;
		color_arr[16167] = 8'b00000000;
		color_arr[16168] = 8'b00000000;
		color_arr[16169] = 8'b00000000;
		color_arr[16170] = 8'b00010010;
		color_arr[16171] = 8'b00010010;
		color_arr[16172] = 8'b00010010;
		color_arr[16173] = 8'b00010010;
		color_arr[16174] = 8'b00010010;
		color_arr[16175] = 8'b00010010;
		color_arr[16176] = 8'b00010010;
		color_arr[16177] = 8'b00010010;
		color_arr[16178] = 8'b00010010;
		color_arr[16179] = 8'b00010010;
		color_arr[16180] = 8'b00010010;
		color_arr[16181] = 8'b00010010;
		color_arr[16182] = 8'b00010010;
		color_arr[16183] = 8'b00010010;
		color_arr[16184] = 8'b00010010;
		color_arr[16185] = 8'b00010010;
		color_arr[16186] = 8'b00010010;
		color_arr[16187] = 8'b00010010;
		color_arr[16188] = 8'b00010010;
		color_arr[16189] = 8'b00010010;
		color_arr[16190] = 8'b00010010;
		color_arr[16191] = 8'b00010010;
		color_arr[16192] = 8'b00010010;
		color_arr[16193] = 8'b00010010;
		color_arr[16194] = 8'b00010010;
		color_arr[16195] = 8'b00010010;
		color_arr[16196] = 8'b00010010;
		color_arr[16197] = 8'b00010010;
		color_arr[16198] = 8'b00010010;
		color_arr[16199] = 8'b00010010;
		color_arr[16200] = 8'b00010010;
		color_arr[16201] = 8'b00010010;
		color_arr[16202] = 8'b00010010;
		color_arr[16203] = 8'b00010010;
		color_arr[16204] = 8'b00010010;
		color_arr[16205] = 8'b00010010;
		color_arr[16206] = 8'b00010010;
		color_arr[16207] = 8'b00010010;
		color_arr[16208] = 8'b00010010;
		color_arr[16209] = 8'b00010010;
		color_arr[16210] = 8'b00010010;
		color_arr[16211] = 8'b00010010;
		color_arr[16212] = 8'b00010010;
		color_arr[16213] = 8'b00010010;
		color_arr[16214] = 8'b00010010;
		color_arr[16215] = 8'b00010010;
		color_arr[16216] = 8'b00010010;
		color_arr[16217] = 8'b00010010;
		color_arr[16218] = 8'b00010010;
		color_arr[16219] = 8'b00010010;
		color_arr[16220] = 8'b00010010;
		color_arr[16221] = 8'b00010010;
		color_arr[16222] = 8'b00010010;
		color_arr[16223] = 8'b00010010;
		color_arr[16224] = 8'b00010010;
		color_arr[16225] = 8'b00010010;
		color_arr[16226] = 8'b00010010;
		color_arr[16227] = 8'b00010010;
		color_arr[16228] = 8'b00010010;
		color_arr[16229] = 8'b00010010;
		color_arr[16230] = 8'b00010010;
		color_arr[16231] = 8'b00010010;
		color_arr[16232] = 8'b00010010;
		color_arr[16233] = 8'b00010010;
		color_arr[16234] = 8'b00010010;
		color_arr[16235] = 8'b00010010;
		color_arr[16236] = 8'b00010010;
		color_arr[16237] = 8'b00010010;
		color_arr[16238] = 8'b00010010;
		color_arr[16239] = 8'b00010010;
		color_arr[16240] = 8'b00010010;
		color_arr[16241] = 8'b00010010;
		color_arr[16242] = 8'b00010010;
		color_arr[16243] = 8'b00010010;
		color_arr[16244] = 8'b00010010;
		color_arr[16245] = 8'b00010010;
		color_arr[16246] = 8'b00010010;
		color_arr[16247] = 8'b00010010;
		color_arr[16248] = 8'b00010010;
		color_arr[16249] = 8'b00010010;
		color_arr[16250] = 8'b00010010;
		color_arr[16251] = 8'b00010010;
		color_arr[16252] = 8'b00010010;
		color_arr[16253] = 8'b00010010;
		color_arr[16254] = 8'b00010010;
		color_arr[16255] = 8'b00010010;
		color_arr[16256] = 8'b00010010;
		color_arr[16257] = 8'b00010010;
		color_arr[16258] = 8'b00010010;
		color_arr[16259] = 8'b00010010;
		color_arr[16260] = 8'b00010010;
		color_arr[16261] = 8'b00010010;
		color_arr[16262] = 8'b00010010;
		color_arr[16263] = 8'b00010010;
		color_arr[16264] = 8'b00010010;
		color_arr[16265] = 8'b00010010;
		color_arr[16266] = 8'b00010010;
		color_arr[16267] = 8'b00010010;
		color_arr[16268] = 8'b00010010;
		color_arr[16269] = 8'b00010010;
		color_arr[16270] = 8'b00010010;
		color_arr[16271] = 8'b00010010;
		color_arr[16272] = 8'b00010010;
		color_arr[16273] = 8'b00010010;
		color_arr[16274] = 8'b00010010;
		color_arr[16275] = 8'b00010010;
		color_arr[16276] = 8'b00010010;
		color_arr[16277] = 8'b00010010;
		color_arr[16278] = 8'b00000000;
		color_arr[16279] = 8'b00000000;
		color_arr[16280] = 8'b00000000;
		color_arr[16281] = 8'b00000000;
		color_arr[16282] = 8'b00000000;
		color_arr[16283] = 8'b00000000;
		color_arr[16284] = 8'b00000000;
		color_arr[16285] = 8'b00000000;
		color_arr[16286] = 8'b00000000;
		color_arr[16287] = 8'b00000000;
		color_arr[16288] = 8'b00000000;
		color_arr[16289] = 8'b00000000;
		color_arr[16290] = 8'b00000000;
		color_arr[16291] = 8'b00000000;
		color_arr[16292] = 8'b00000000;
		color_arr[16293] = 8'b00000000;
		color_arr[16294] = 8'b00000000;
		color_arr[16295] = 8'b00000000;
		color_arr[16296] = 8'b00010010;
		color_arr[16297] = 8'b00010010;
		color_arr[16298] = 8'b00010010;
		color_arr[16299] = 8'b00010010;
		color_arr[16300] = 8'b00010010;
		color_arr[16301] = 8'b00010010;
		color_arr[16302] = 8'b00010010;
		color_arr[16303] = 8'b00010010;
		color_arr[16304] = 8'b00010010;
		color_arr[16305] = 8'b00010010;
		color_arr[16306] = 8'b00010010;
		color_arr[16307] = 8'b00010010;
		color_arr[16308] = 8'b00010010;
		color_arr[16309] = 8'b00010010;
		color_arr[16310] = 8'b00010010;
		color_arr[16311] = 8'b00010010;
		color_arr[16312] = 8'b00010010;
		color_arr[16313] = 8'b00010010;
		color_arr[16314] = 8'b00010010;
		color_arr[16315] = 8'b00010010;
		color_arr[16316] = 8'b00010010;
		color_arr[16317] = 8'b00010010;
		color_arr[16318] = 8'b00010010;
		color_arr[16319] = 8'b00010010;
		color_arr[16320] = 8'b00010010;
		color_arr[16321] = 8'b00010010;
		color_arr[16322] = 8'b00010010;
		color_arr[16323] = 8'b00010010;
		color_arr[16324] = 8'b00010010;
		color_arr[16325] = 8'b00010010;
		color_arr[16326] = 8'b00010010;
		color_arr[16327] = 8'b00010010;
		color_arr[16328] = 8'b00010010;
		color_arr[16329] = 8'b00010010;
		color_arr[16330] = 8'b00010010;
		color_arr[16331] = 8'b00010010;
		color_arr[16332] = 8'b00010010;
		color_arr[16333] = 8'b00010010;
		color_arr[16334] = 8'b00010010;
		color_arr[16335] = 8'b00010010;
		color_arr[16336] = 8'b00010010;
		color_arr[16337] = 8'b00010010;
		color_arr[16338] = 8'b00010010;
		color_arr[16339] = 8'b00010010;
		color_arr[16340] = 8'b00010010;
		color_arr[16341] = 8'b00010010;
		color_arr[16342] = 8'b00010010;
		color_arr[16343] = 8'b00010010;
		color_arr[16344] = 8'b00010010;
		color_arr[16345] = 8'b00010010;
		color_arr[16346] = 8'b00010010;
		color_arr[16347] = 8'b00010010;
		color_arr[16348] = 8'b00010010;
		color_arr[16349] = 8'b00010010;
		color_arr[16350] = 8'b00010010;
		color_arr[16351] = 8'b00010010;
		color_arr[16352] = 8'b00010010;
		color_arr[16353] = 8'b00010010;
		color_arr[16354] = 8'b00010010;
		color_arr[16355] = 8'b00010010;
		color_arr[16356] = 8'b00010010;
		color_arr[16357] = 8'b00010010;
		color_arr[16358] = 8'b00010010;
		color_arr[16359] = 8'b00010010;
		color_arr[16360] = 8'b00010010;
		color_arr[16361] = 8'b00010010;
		color_arr[16362] = 8'b00010010;
		color_arr[16363] = 8'b00010010;
		color_arr[16364] = 8'b00010010;
		color_arr[16365] = 8'b00010010;
		color_arr[16366] = 8'b00010010;
		color_arr[16367] = 8'b00010010;
		color_arr[16368] = 8'b00010010;
		color_arr[16369] = 8'b00010010;
		color_arr[16370] = 8'b00010010;
		color_arr[16371] = 8'b00010010;
		color_arr[16372] = 8'b00010010;
		color_arr[16373] = 8'b00010010;
		color_arr[16374] = 8'b00010010;
		color_arr[16375] = 8'b00010010;
		color_arr[16376] = 8'b00010010;
		color_arr[16377] = 8'b00010010;
		color_arr[16378] = 8'b00010010;
		color_arr[16379] = 8'b00010010;
		color_arr[16380] = 8'b00010010;
		color_arr[16381] = 8'b00010010;
		color_arr[16382] = 8'b00010010;
		color_arr[16383] = 8'b00010010;
	end

	always @(posedge clk) begin
		color_out <= color_arr[addr][5:0];
	end
endmodule
